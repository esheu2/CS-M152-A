`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    09:41:20 03/07/2019 
// Design Name: 
// Module Name:    sigmoid_approx 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
// Implemented sigmoid with piece-wise linear approximation from http://www.iosrjen.org/Papers/vol2_issue6%20(part-1)/N026135521356.pdf
// This is much easier for the FPGA to compute
module sigmoid_approx(
	clk,
	x,
	y);

input clk;	
	
input wire [31:0] x;
output wire [31:0] y;

reg [31:0] y_temp;

always@(x)
begin
if(x[31] == 0)
begin
if( x > 32'b00000000000000000000000000000000 && x < 32'b00111100001000111101011100001010)
begin
	y_temp <= 32'b00111111000000000101000111101011;
end
if( x >= 32'b00111100001000111101011100001010 && x < 32'b00111100101000111101011100001010)
begin
	y_temp <= 32'b00111111000000001111010111000001;
end
if( x >= 32'b00111100101000111101011100001010 && x < 32'b00111100111101011100001010001111)
begin
	y_temp <= 32'b00111111000000011001100110010100;
end
if( x >= 32'b00111100111101011100001010001111 && x < 32'b00111101001000111101011100001010)
begin
	y_temp <= 32'b00111111000000100011110101100010;
end
if( x >= 32'b00111101001000111101011100001010 && x < 32'b00111101010011001100110011001101)
begin
	y_temp <= 32'b00111111000000101110000100101000;
end
if( x >= 32'b00111101010011001100110011001101 && x < 32'b00111101011101011100001010001111)
begin
	y_temp <= 32'b00111111000000111000010011100101;
end
if( x >= 32'b00111101011101011100001010001111 && x < 32'b00111101100011110101110000101001)
begin
	y_temp <= 32'b00111111000001000010100010010110;
end
if( x >= 32'b00111101100011110101110000101001 && x < 32'b00111101101000111101011100001010)
begin
	y_temp <= 32'b00111111000001001100110000111001;
end
if( x >= 32'b00111101101000111101011100001010 && x < 32'b00111101101110000101000111101100)
begin
	y_temp <= 32'b00111111000001010110111111001101;
end
if( x >= 32'b00111101101110000101000111101100 && x < 32'b00111101110011001100110011001101)
begin
	y_temp <= 32'b00111111000001100001001101001111;
end
if( x >= 32'b00111101110011001100110011001101 && x < 32'b00111101111000010100011110101110)
begin
	y_temp <= 32'b00111111000001101011011010111110;
end
if( x >= 32'b00111101111000010100011110101110 && x < 32'b00111101111101011100001010001111)
begin
	y_temp <= 32'b00111111000001110101101000010110;
end
if( x >= 32'b00111101111101011100001010001111 && x < 32'b00111110000001010001111010111000)
begin
	y_temp <= 32'b00111111000001111111110101010110;
end
if( x >= 32'b00111110000001010001111010111000 && x < 32'b00111110000011110101110000101001)
begin
	y_temp <= 32'b00111111000010001010000001111101;
end
if( x >= 32'b00111110000011110101110000101001 && x < 32'b00111110000110011001100110011010)
begin
	y_temp <= 32'b00111111000010010100001110000111;
end
if( x >= 32'b00111110000110011001100110011010 && x < 32'b00111110001000111101011100001010)
begin
	y_temp <= 32'b00111111000010011110011001110011;
end
if( x >= 32'b00111110001000111101011100001010 && x < 32'b00111110001011100001010001111011)
begin
	y_temp <= 32'b00111111000010101000100100111110;
end
if( x >= 32'b00111110001011100001010001111011 && x < 32'b00111110001110000101000111101100)
begin
	y_temp <= 32'b00111111000010110010101111101000;
end
if( x >= 32'b00111110001110000101000111101100 && x < 32'b00111110010000101000111101011100)
begin
	y_temp <= 32'b00111111000010111100111001101101;
end
if( x >= 32'b00111110010000101000111101011100 && x < 32'b00111110010011001100110011001101)
begin
	y_temp <= 32'b00111111000011000111000011001011;
end
if( x >= 32'b00111110010011001100110011001101 && x < 32'b00111110010101110000101000111101)
begin
	y_temp <= 32'b00111111000011010001001100000010;
end
if( x >= 32'b00111110010101110000101000111101 && x < 32'b00111110011000010100011110101110)
begin
	y_temp <= 32'b00111111000011011011010100001110;
end
if( x >= 32'b00111110011000010100011110101110 && x < 32'b00111110011010111000010100011111)
begin
	y_temp <= 32'b00111111000011100101011011101101;
end
if( x >= 32'b00111110011010111000010100011111 && x < 32'b00111110011101011100001010001111)
begin
	y_temp <= 32'b00111111000011101111100010011110;
end
if( x >= 32'b00111110011101011100001010001111 && x < 32'b00111110100000000000000000000000)
begin
	y_temp <= 32'b00111111000011111001101000011111;
end
if( x >= 32'b00111110100000000000000000000000 && x < 32'b00111110100001010001111010111000)
begin
	y_temp <= 32'b00111111000100000011101101101101;
end
if( x >= 32'b00111110100001010001111010111000 && x < 32'b00111110100010100011110101110001)
begin
	y_temp <= 32'b00111111000100001101110010000111;
end
if( x >= 32'b00111110100010100011110101110001 && x < 32'b00111110100011110101110000101001)
begin
	y_temp <= 32'b00111111000100010111110101101011;
end
if( x >= 32'b00111110100011110101110000101001 && x < 32'b00111110100101000111101011100001)
begin
	y_temp <= 32'b00111111000100100001111000010111;
end
if( x >= 32'b00111110100101000111101011100001 && x < 32'b00111110100110011001100110011010)
begin
	y_temp <= 32'b00111111000100101011111010001000;
end
if( x >= 32'b00111110100110011001100110011010 && x < 32'b00111110100111101011100001010010)
begin
	y_temp <= 32'b00111111000100110101111010111101;
end
if( x >= 32'b00111110100111101011100001010010 && x < 32'b00111110101000111101011100001010)
begin
	y_temp <= 32'b00111111000100111111111010110100;
end
if( x >= 32'b00111110101000111101011100001010 && x < 32'b00111110101010001111010111000011)
begin
	y_temp <= 32'b00111111000101001001111001101100;
end
if( x >= 32'b00111110101010001111010111000011 && x < 32'b00111110101011100001010001111011)
begin
	y_temp <= 32'b00111111000101010011110111100001;
end
if( x >= 32'b00111110101011100001010001111011 && x < 32'b00111110101100110011001100110011)
begin
	y_temp <= 32'b00111111000101011101110100010011;
end
if( x >= 32'b00111110101100110011001100110011 && x < 32'b00111110101110000101000111101100)
begin
	y_temp <= 32'b00111111000101100111101111111111;
end
if( x >= 32'b00111110101110000101000111101100 && x < 32'b00111110101111010111000010100100)
begin
	y_temp <= 32'b00111111000101110001101010100100;
end
if( x >= 32'b00111110101111010111000010100100 && x < 32'b00111110110000101000111101011100)
begin
	y_temp <= 32'b00111111000101111011100100000000;
end
if( x >= 32'b00111110110000101000111101011100 && x < 32'b00111110110001111010111000010100)
begin
	y_temp <= 32'b00111111000110000101011100010000;
end
if( x >= 32'b00111110110001111010111000010100 && x < 32'b00111110110011001100110011001101)
begin
	y_temp <= 32'b00111111000110001111010011010100;
end
if( x >= 32'b00111110110011001100110011001101 && x < 32'b00111110110100011110101110000101)
begin
	y_temp <= 32'b00111111000110011001001001001001;
end
if( x >= 32'b00111110110100011110101110000101 && x < 32'b00111110110101110000101000111101)
begin
	y_temp <= 32'b00111111000110100010111101101101;
end
if( x >= 32'b00111110110101110000101000111101 && x < 32'b00111110110111000010100011110110)
begin
	y_temp <= 32'b00111111000110101100110001000000;
end
if( x >= 32'b00111110110111000010100011110110 && x < 32'b00111110111000010100011110101110)
begin
	y_temp <= 32'b00111111000110110110100010111110;
end
if( x >= 32'b00111110111000010100011110101110 && x < 32'b00111110111001100110011001100110)
begin
	y_temp <= 32'b00111111000111000000010011100111;
end
if( x >= 32'b00111110111001100110011001100110 && x < 32'b00111110111010111000010100011111)
begin
	y_temp <= 32'b00111111000111001010000010111000;
end
if( x >= 32'b00111110111010111000010100011111 && x < 32'b00111110111100001010001111010111)
begin
	y_temp <= 32'b00111111000111010011110000110000;
end
if( x >= 32'b00111110111100001010001111010111 && x < 32'b00111110111101011100001010001111)
begin
	y_temp <= 32'b00111111000111011101011101001101;
end
if( x >= 32'b00111110111101011100001010001111 && x < 32'b00111110111110101110000101001000)
begin
	y_temp <= 32'b00111111000111100111001000001110;
end
if( x >= 32'b00111110111110101110000101001000 && x < 32'b00111111000000000000000000000000)
begin
	y_temp <= 32'b00111111000111110000110001110001;
end
if( x >= 32'b00111111000000000000000000000000 && x < 32'b00111111000000101000111101011100)
begin
	y_temp <= 32'b00111111000111111010011001110100;
end
if( x >= 32'b00111111000000101000111101011100 && x < 32'b00111111000001010001111010111000)
begin
	y_temp <= 32'b00111111001000000100000000010110;
end
if( x >= 32'b00111111000001010001111010111000 && x < 32'b00111111000001111010111000010100)
begin
	y_temp <= 32'b00111111001000001101100101010100;
end
if( x >= 32'b00111111000001111010111000010100 && x < 32'b00111111000010100011110101110001)
begin
	y_temp <= 32'b00111111001000010111001000101111;
end
if( x >= 32'b00111111000010100011110101110001 && x < 32'b00111111000011001100110011001101)
begin
	y_temp <= 32'b00111111001000100000101010100011;
end
if( x >= 32'b00111111000011001100110011001101 && x < 32'b00111111000011110101110000101001)
begin
	y_temp <= 32'b00111111001000101010001010101111;
end
if( x >= 32'b00111111000011110101110000101001 && x < 32'b00111111000100011110101110000101)
begin
	y_temp <= 32'b00111111001000110011101001010010;
end
if( x >= 32'b00111111000100011110101110000101 && x < 32'b00111111000101000111101011100001)
begin
	y_temp <= 32'b00111111001000111101000110001011;
end
if( x >= 32'b00111111000101000111101011100001 && x < 32'b00111111000101110000101000111101)
begin
	y_temp <= 32'b00111111001001000110100001010111;
end
if( x >= 32'b00111111000101110000101000111101 && x < 32'b00111111000110011001100110011010)
begin
	y_temp <= 32'b00111111001001001111111010110110;
end
if( x >= 32'b00111111000110011001100110011010 && x < 32'b00111111000111000010100011110110)
begin
	y_temp <= 32'b00111111001001011001010010100101;
end
if( x >= 32'b00111111000111000010100011110110 && x < 32'b00111111000111101011100001010010)
begin
	y_temp <= 32'b00111111001001100010101000100100;
end
if( x >= 32'b00111111000111101011100001010010 && x < 32'b00111111001000010100011110101110)
begin
	y_temp <= 32'b00111111001001101011111100110001;
end
if( x >= 32'b00111111001000010100011110101110 && x < 32'b00111111001000111101011100001010)
begin
	y_temp <= 32'b00111111001001110101001111001011;
end
if( x >= 32'b00111111001000111101011100001010 && x < 32'b00111111001001100110011001100110)
begin
	y_temp <= 32'b00111111001001111110011111110000;
end
if( x >= 32'b00111111001001100110011001100110 && x < 32'b00111111001010001111010111000011)
begin
	y_temp <= 32'b00111111001010000111101110011111;
end
if( x >= 32'b00111111001010001111010111000011 && x < 32'b00111111001010111000010100011111)
begin
	y_temp <= 32'b00111111001010010000111011010111;
end
if( x >= 32'b00111111001010111000010100011111 && x < 32'b00111111001011100001010001111011)
begin
	y_temp <= 32'b00111111001010011010000110010110;
end
if( x >= 32'b00111111001011100001010001111011 && x < 32'b00111111001100001010001111010111)
begin
	y_temp <= 32'b00111111001010100011001111011011;
end
if( x >= 32'b00111111001100001010001111010111 && x < 32'b00111111001100110011001100110011)
begin
	y_temp <= 32'b00111111001010101100010110100100;
end
if( x >= 32'b00111111001100110011001100110011 && x < 32'b00111111001101011100001010001111)
begin
	y_temp <= 32'b00111111001010110101011011110010;
end
if( x >= 32'b00111111001101011100001010001111 && x < 32'b00111111001110000101000111101100)
begin
	y_temp <= 32'b00111111001010111110011111000001;
end
if( x >= 32'b00111111001110000101000111101100 && x < 32'b00111111001110101110000101001000)
begin
	y_temp <= 32'b00111111001011000111100000010010;
end
if( x >= 32'b00111111001110101110000101001000 && x < 32'b00111111001111010111000010100100)
begin
	y_temp <= 32'b00111111001011010000011111100010;
end
if( x >= 32'b00111111001111010111000010100100 && x < 32'b00111111010000000000000000000000)
begin
	y_temp <= 32'b00111111001011011001011100110001;
end
if( x >= 32'b00111111010000000000000000000000 && x < 32'b00111111010000101000111101011100)
begin
	y_temp <= 32'b00111111001011100010010111111110;
end
if( x >= 32'b00111111010000101000111101011100 && x < 32'b00111111010001010001111010111000)
begin
	y_temp <= 32'b00111111001011101011010001000111;
end
if( x >= 32'b00111111010001010001111010111000 && x < 32'b00111111010001111010111000010100)
begin
	y_temp <= 32'b00111111001011110100001000001011;
end
if( x >= 32'b00111111010001111010111000010100 && x < 32'b00111111010010100011110101110001)
begin
	y_temp <= 32'b00111111001011111100111101001010;
end
if( x >= 32'b00111111010010100011110101110001 && x < 32'b00111111010011001100110011001101)
begin
	y_temp <= 32'b00111111001100000101110000000010;
end
if( x >= 32'b00111111010011001100110011001101 && x < 32'b00111111010011110101110000101001)
begin
	y_temp <= 32'b00111111001100001110100000110010;
end
if( x >= 32'b00111111010011110101110000101001 && x < 32'b00111111010100011110101110000101)
begin
	y_temp <= 32'b00111111001100010111001111011001;
end
if( x >= 32'b00111111010100011110101110000101 && x < 32'b00111111010101000111101011100001)
begin
	y_temp <= 32'b00111111001100011111111011110110;
end
if( x >= 32'b00111111010101000111101011100001 && x < 32'b00111111010101110000101000111101)
begin
	y_temp <= 32'b00111111001100101000100110001001;
end
if( x >= 32'b00111111010101110000101000111101 && x < 32'b00111111010110011001100110011010)
begin
	y_temp <= 32'b00111111001100110001001110010000;
end
if( x >= 32'b00111111010110011001100110011010 && x < 32'b00111111010111000010100011110110)
begin
	y_temp <= 32'b00111111001100111001110100001010;
end
if( x >= 32'b00111111010111000010100011110110 && x < 32'b00111111010111101011100001010010)
begin
	y_temp <= 32'b00111111001101000010010111110110;
end
if( x >= 32'b00111111010111101011100001010010 && x < 32'b00111111011000010100011110101110)
begin
	y_temp <= 32'b00111111001101001010111001010100;
end
if( x >= 32'b00111111011000010100011110101110 && x < 32'b00111111011000111101011100001010)
begin
	y_temp <= 32'b00111111001101010011011000100010;
end
if( x >= 32'b00111111011000111101011100001010 && x < 32'b00111111011001100110011001100110)
begin
	y_temp <= 32'b00111111001101011011110101100001;
end
if( x >= 32'b00111111011001100110011001100110 && x < 32'b00111111011010001111010111000011)
begin
	y_temp <= 32'b00111111001101100100010000001110;
end
if( x >= 32'b00111111011010001111010111000011 && x < 32'b00111111011010111000010100011111)
begin
	y_temp <= 32'b00111111001101101100101000101001;
end
if( x >= 32'b00111111011010111000010100011111 && x < 32'b00111111011011100001010001111011)
begin
	y_temp <= 32'b00111111001101110100111110110010;
end
if( x >= 32'b00111111011011100001010001111011 && x < 32'b00111111011100001010001111010111)
begin
	y_temp <= 32'b00111111001101111101010010100111;
end
if( x >= 32'b00111111011100001010001111010111 && x < 32'b00111111011100110011001100110011)
begin
	y_temp <= 32'b00111111001110000101100100001000;
end
if( x >= 32'b00111111011100110011001100110011 && x < 32'b00111111011101011100001010001111)
begin
	y_temp <= 32'b00111111001110001101110011010101;
end
if( x >= 32'b00111111011101011100001010001111 && x < 32'b00111111011110000101000111101100)
begin
	y_temp <= 32'b00111111001110010110000000001011;
end
if( x >= 32'b00111111011110000101000111101100 && x < 32'b00111111011110101110000101001000)
begin
	y_temp <= 32'b00111111001110011110001010101100;
end
if( x >= 32'b00111111011110101110000101001000 && x < 32'b00111111011111010111000010100100)
begin
	y_temp <= 32'b00111111001110100110010010110110;
end
if( x >= 32'b00111111011111010111000010100100 && x < 32'b00111111100000000000000000000000)
begin
	y_temp <= 32'b00111111001110101110011000101000;
end
if( x >= 32'b00111111100000000000000000000000 && x < 32'b00111111100000010100011110101110)
begin
	y_temp <= 32'b00111111001110110110011100000010;
end
if( x >= 32'b00111111100000010100011110101110 && x < 32'b00111111100000101000111101011100)
begin
	y_temp <= 32'b00111111001110111110011101000011;
end
if( x >= 32'b00111111100000101000111101011100 && x < 32'b00111111100000111101011100001010)
begin
	y_temp <= 32'b00111111001111000110011011101011;
end
if( x >= 32'b00111111100000111101011100001010 && x < 32'b00111111100001010001111010111000)
begin
	y_temp <= 32'b00111111001111001110010111111001;
end
if( x >= 32'b00111111100001010001111010111000 && x < 32'b00111111100001100110011001100110)
begin
	y_temp <= 32'b00111111001111010110010001101101;
end
if( x >= 32'b00111111100001100110011001100110 && x < 32'b00111111100001111010111000010100)
begin
	y_temp <= 32'b00111111001111011110001001000110;
end
if( x >= 32'b00111111100001111010111000010100 && x < 32'b00111111100010001111010111000011)
begin
	y_temp <= 32'b00111111001111100101111110000011;
end
if( x >= 32'b00111111100010001111010111000011 && x < 32'b00111111100010100011110101110001)
begin
	y_temp <= 32'b00111111001111101101110000100101;
end
if( x >= 32'b00111111100010100011110101110001 && x < 32'b00111111100010111000010100011111)
begin
	y_temp <= 32'b00111111001111110101100000101010;
end
if( x >= 32'b00111111100010111000010100011111 && x < 32'b00111111100011001100110011001101)
begin
	y_temp <= 32'b00111111001111111101001110010010;
end
if( x >= 32'b00111111100011001100110011001101 && x < 32'b00111111100011100001010001111011)
begin
	y_temp <= 32'b00111111010000000100111001011110;
end
if( x >= 32'b00111111100011100001010001111011 && x < 32'b00111111100011110101110000101001)
begin
	y_temp <= 32'b00111111010000001100100010001100;
end
if( x >= 32'b00111111100011110101110000101001 && x < 32'b00111111100100001010001111010111)
begin
	y_temp <= 32'b00111111010000010100001000011100;
end
if( x >= 32'b00111111100100001010001111010111 && x < 32'b00111111100100011110101110000101)
begin
	y_temp <= 32'b00111111010000011011101100001110;
end
if( x >= 32'b00111111100100011110101110000101 && x < 32'b00111111100100110011001100110011)
begin
	y_temp <= 32'b00111111010000100011001101100001;
end
if( x >= 32'b00111111100100110011001100110011 && x < 32'b00111111100101000111101011100001)
begin
	y_temp <= 32'b00111111010000101010101100010101;
end
if( x >= 32'b00111111100101000111101011100001 && x < 32'b00111111100101011100001010001111)
begin
	y_temp <= 32'b00111111010000110010001000101010;
end
if( x >= 32'b00111111100101011100001010001111 && x < 32'b00111111100101110000101000111101)
begin
	y_temp <= 32'b00111111010000111001100010100000;
end
if( x >= 32'b00111111100101110000101000111101 && x < 32'b00111111100110000101000111101100)
begin
	y_temp <= 32'b00111111010001000000111001110101;
end
if( x >= 32'b00111111100110000101000111101100 && x < 32'b00111111100110011001100110011010)
begin
	y_temp <= 32'b00111111010001001000001110101011;
end
if( x >= 32'b00111111100110011001100110011010 && x < 32'b00111111100110101110000101001000)
begin
	y_temp <= 32'b00111111010001001111100001000001;
end
if( x >= 32'b00111111100110101110000101001000 && x < 32'b00111111100111000010100011110110)
begin
	y_temp <= 32'b00111111010001010110110000110110;
end
if( x >= 32'b00111111100111000010100011110110 && x < 32'b00111111100111010111000010100100)
begin
	y_temp <= 32'b00111111010001011101111110001011;
end
if( x >= 32'b00111111100111010111000010100100 && x < 32'b00111111100111101011100001010010)
begin
	y_temp <= 32'b00111111010001100101001000111111;
end
if( x >= 32'b00111111100111101011100001010010 && x < 32'b00111111101000000000000000000000)
begin
	y_temp <= 32'b00111111010001101100010001010010;
end
if( x >= 32'b00111111101000000000000000000000 && x < 32'b00111111101000010100011110101110)
begin
	y_temp <= 32'b00111111010001110011010111000101;
end
if( x >= 32'b00111111101000010100011110101110 && x < 32'b00111111101000101000111101011100)
begin
	y_temp <= 32'b00111111010001111010011010010110;
end
if( x >= 32'b00111111101000101000111101011100 && x < 32'b00111111101000111101011100001010)
begin
	y_temp <= 32'b00111111010010000001011011000101;
end
if( x >= 32'b00111111101000111101011100001010 && x < 32'b00111111101001010001111010111000)
begin
	y_temp <= 32'b00111111010010001000011001010100;
end
if( x >= 32'b00111111101001010001111010111000 && x < 32'b00111111101001100110011001100110)
begin
	y_temp <= 32'b00111111010010001111010101000001;
end
if( x >= 32'b00111111101001100110011001100110 && x < 32'b00111111101001111010111000010100)
begin
	y_temp <= 32'b00111111010010010110001110001101;
end
if( x >= 32'b00111111101001111010111000010100 && x < 32'b00111111101010001111010111000011)
begin
	y_temp <= 32'b00111111010010011101000100110111;
end
if( x >= 32'b00111111101010001111010111000011 && x < 32'b00111111101010100011110101110001)
begin
	y_temp <= 32'b00111111010010100011111001000000;
end
if( x >= 32'b00111111101010100011110101110001 && x < 32'b00111111101010111000010100011111)
begin
	y_temp <= 32'b00111111010010101010101010101000;
end
if( x >= 32'b00111111101010111000010100011111 && x < 32'b00111111101011001100110011001101)
begin
	y_temp <= 32'b00111111010010110001011001101110;
end
if( x >= 32'b00111111101011001100110011001101 && x < 32'b00111111101011100001010001111011)
begin
	y_temp <= 32'b00111111010010111000000110010010;
end
if( x >= 32'b00111111101011100001010001111011 && x < 32'b00111111101011110101110000101001)
begin
	y_temp <= 32'b00111111010010111110110000010110;
end
if( x >= 32'b00111111101011110101110000101001 && x < 32'b00111111101100001010001111010111)
begin
	y_temp <= 32'b00111111010011000101010111111000;
end
if( x >= 32'b00111111101100001010001111010111 && x < 32'b00111111101100011110101110000101)
begin
	y_temp <= 32'b00111111010011001011111100111001;
end
if( x >= 32'b00111111101100011110101110000101 && x < 32'b00111111101100110011001100110011)
begin
	y_temp <= 32'b00111111010011010010011111011001;
end
if( x >= 32'b00111111101100110011001100110011 && x < 32'b00111111101101000111101011100001)
begin
	y_temp <= 32'b00111111010011011000111111011000;
end
if( x >= 32'b00111111101101000111101011100001 && x < 32'b00111111101101011100001010001111)
begin
	y_temp <= 32'b00111111010011011111011100110110;
end
if( x >= 32'b00111111101101011100001010001111 && x < 32'b00111111101101110000101000111101)
begin
	y_temp <= 32'b00111111010011100101110111110011;
end
if( x >= 32'b00111111101101110000101000111101 && x < 32'b00111111101110000101000111101100)
begin
	y_temp <= 32'b00111111010011101100010000010000;
end
if( x >= 32'b00111111101110000101000111101100 && x < 32'b00111111101110011001100110011010)
begin
	y_temp <= 32'b00111111010011110010100110001101;
end
if( x >= 32'b00111111101110011001100110011010 && x < 32'b00111111101110101110000101001000)
begin
	y_temp <= 32'b00111111010011111000111001101001;
end
if( x >= 32'b00111111101110101110000101001000 && x < 32'b00111111101111000010100011110110)
begin
	y_temp <= 32'b00111111010011111111001010100101;
end
if( x >= 32'b00111111101111000010100011110110 && x < 32'b00111111101111010111000010100100)
begin
	y_temp <= 32'b00111111010100000101011001000010;
end
if( x >= 32'b00111111101111010111000010100100 && x < 32'b00111111101111101011100001010010)
begin
	y_temp <= 32'b00111111010100001011100100111111;
end
if( x >= 32'b00111111101111101011100001010010 && x < 32'b00111111110000000000000000000000)
begin
	y_temp <= 32'b00111111010100010001101110011100;
end
if( x >= 32'b00111111110000000000000000000000 && x < 32'b00111111110000010100011110101110)
begin
	y_temp <= 32'b00111111010100010111110101011011;
end
if( x >= 32'b00111111110000010100011110101110 && x < 32'b00111111110000101000111101011100)
begin
	y_temp <= 32'b00111111010100011101111001111011;
end
if( x >= 32'b00111111110000101000111101011100 && x < 32'b00111111110000111101011100001010)
begin
	y_temp <= 32'b00111111010100100011111011111100;
end
if( x >= 32'b00111111110000111101011100001010 && x < 32'b00111111110001010001111010111000)
begin
	y_temp <= 32'b00111111010100101001111011011111;
end
if( x >= 32'b00111111110001010001111010111000 && x < 32'b00111111110001100110011001100110)
begin
	y_temp <= 32'b00111111010100101111111000100100;
end
if( x >= 32'b00111111110001100110011001100110 && x < 32'b00111111110001111010111000010100)
begin
	y_temp <= 32'b00111111010100110101110011001100;
end
if( x >= 32'b00111111110001111010111000010100 && x < 32'b00111111110010001111010111000011)
begin
	y_temp <= 32'b00111111010100111011101011010110;
end
if( x >= 32'b00111111110010001111010111000011 && x < 32'b00111111110010100011110101110001)
begin
	y_temp <= 32'b00111111010101000001100001000011;
end
if( x >= 32'b00111111110010100011110101110001 && x < 32'b00111111110010111000010100011111)
begin
	y_temp <= 32'b00111111010101000111010100010100;
end
if( x >= 32'b00111111110010111000010100011111 && x < 32'b00111111110011001100110011001101)
begin
	y_temp <= 32'b00111111010101001101000101001000;
end
if( x >= 32'b00111111110011001100110011001101 && x < 32'b00111111110011100001010001111011)
begin
	y_temp <= 32'b00111111010101010010110011100001;
end
if( x >= 32'b00111111110011100001010001111011 && x < 32'b00111111110011110101110000101001)
begin
	y_temp <= 32'b00111111010101011000011111011110;
end
if( x >= 32'b00111111110011110101110000101001 && x < 32'b00111111110100001010001111010111)
begin
	y_temp <= 32'b00111111010101011110001001000000;
end
if( x >= 32'b00111111110100001010001111010111 && x < 32'b00111111110100011110101110000101)
begin
	y_temp <= 32'b00111111010101100011110000000111;
end
if( x >= 32'b00111111110100011110101110000101 && x < 32'b00111111110100110011001100110011)
begin
	y_temp <= 32'b00111111010101101001010100110100;
end
if( x >= 32'b00111111110100110011001100110011 && x < 32'b00111111110101000111101011100001)
begin
	y_temp <= 32'b00111111010101101110110111000111;
end
if( x >= 32'b00111111110101000111101011100001 && x < 32'b00111111110101011100001010001111)
begin
	y_temp <= 32'b00111111010101110100010111000000;
end
if( x >= 32'b00111111110101011100001010001111 && x < 32'b00111111110101110000101000111101)
begin
	y_temp <= 32'b00111111010101111001110100100000;
end
if( x >= 32'b00111111110101110000101000111101 && x < 32'b00111111110110000101000111101100)
begin
	y_temp <= 32'b00111111010101111111001111101000;
end
if( x >= 32'b00111111110110000101000111101100 && x < 32'b00111111110110011001100110011010)
begin
	y_temp <= 32'b00111111010110000100101000011000;
end
if( x >= 32'b00111111110110011001100110011010 && x < 32'b00111111110110101110000101001000)
begin
	y_temp <= 32'b00111111010110001001111110110000;
end
if( x >= 32'b00111111110110101110000101001000 && x < 32'b00111111110111000010100011110110)
begin
	y_temp <= 32'b00111111010110001111010010110001;
end
if( x >= 32'b00111111110111000010100011110110 && x < 32'b00111111110111010111000010100100)
begin
	y_temp <= 32'b00111111010110010100100100011011;
end
if( x >= 32'b00111111110111010111000010100100 && x < 32'b00111111110111101011100001010010)
begin
	y_temp <= 32'b00111111010110011001110011101111;
end
if( x >= 32'b00111111110111101011100001010010 && x < 32'b00111111111000000000000000000000)
begin
	y_temp <= 32'b00111111010110011111000000101101;
end
if( x >= 32'b00111111111000000000000000000000 && x < 32'b00111111111000010100011110101110)
begin
	y_temp <= 32'b00111111010110100100001011010110;
end
if( x >= 32'b00111111111000010100011110101110 && x < 32'b00111111111000101000111101011100)
begin
	y_temp <= 32'b00111111010110101001010011101010;
end
if( x >= 32'b00111111111000101000111101011100 && x < 32'b00111111111000111101011100001010)
begin
	y_temp <= 32'b00111111010110101110011001101010;
end
if( x >= 32'b00111111111000111101011100001010 && x < 32'b00111111111001010001111010111000)
begin
	y_temp <= 32'b00111111010110110011011101010111;
end
if( x >= 32'b00111111111001010001111010111000 && x < 32'b00111111111001100110011001100110)
begin
	y_temp <= 32'b00111111010110111000011110110000;
end
if( x >= 32'b00111111111001100110011001100110 && x < 32'b00111111111001111010111000010100)
begin
	y_temp <= 32'b00111111010110111101011101110111;
end
if( x >= 32'b00111111111001111010111000010100 && x < 32'b00111111111010001111010111000011)
begin
	y_temp <= 32'b00111111010111000010011010101100;
end
if( x >= 32'b00111111111010001111010111000011 && x < 32'b00111111111010100011110101110001)
begin
	y_temp <= 32'b00111111010111000111010101001111;
end
if( x >= 32'b00111111111010100011110101110001 && x < 32'b00111111111010111000010100011111)
begin
	y_temp <= 32'b00111111010111001100001101100010;
end
if( x >= 32'b00111111111010111000010100011111 && x < 32'b00111111111011001100110011001101)
begin
	y_temp <= 32'b00111111010111010001000011100100;
end
if( x >= 32'b00111111111011001100110011001101 && x < 32'b00111111111011100001010001111011)
begin
	y_temp <= 32'b00111111010111010101110111010110;
end
if( x >= 32'b00111111111011100001010001111011 && x < 32'b00111111111011110101110000101001)
begin
	y_temp <= 32'b00111111010111011010101000111010;
end
if( x >= 32'b00111111111011110101110000101001 && x < 32'b00111111111100001010001111010111)
begin
	y_temp <= 32'b00111111010111011111011000001110;
end
if( x >= 32'b00111111111100001010001111010111 && x < 32'b00111111111100011110101110000101)
begin
	y_temp <= 32'b00111111010111100100000101010101;
end
if( x >= 32'b00111111111100011110101110000101 && x < 32'b00111111111100110011001100110011)
begin
	y_temp <= 32'b00111111010111101000110000001110;
end
if( x >= 32'b00111111111100110011001100110011 && x < 32'b00111111111101000111101011100001)
begin
	y_temp <= 32'b00111111010111101101011000111011;
end
if( x >= 32'b00111111111101000111101011100001 && x < 32'b00111111111101011100001010001111)
begin
	y_temp <= 32'b00111111010111110001111111011011;
end
if( x >= 32'b00111111111101011100001010001111 && x < 32'b00111111111101110000101000111101)
begin
	y_temp <= 32'b00111111010111110110100011110000;
end
if( x >= 32'b00111111111101110000101000111101 && x < 32'b00111111111110000101000111101100)
begin
	y_temp <= 32'b00111111010111111011000101111010;
end
if( x >= 32'b00111111111110000101000111101100 && x < 32'b00111111111110011001100110011010)
begin
	y_temp <= 32'b00111111010111111111100101111001;
end
if( x >= 32'b00111111111110011001100110011010 && x < 32'b00111111111110101110000101001000)
begin
	y_temp <= 32'b00111111011000000100000011101111;
end
if( x >= 32'b00111111111110101110000101001000 && x < 32'b00111111111111000010100011110110)
begin
	y_temp <= 32'b00111111011000001000011111011100;
end
if( x >= 32'b00111111111111000010100011110110 && x < 32'b00111111111111010111000010100100)
begin
	y_temp <= 32'b00111111011000001100111001000000;
end
if( x >= 32'b00111111111111010111000010100100 && x < 32'b00111111111111101011100001010010)
begin
	y_temp <= 32'b00111111011000010001010000011101;
end
if( x >= 32'b00111111111111101011100001010010 && x < 32'b01000000000000000000000000000000)
begin
	y_temp <= 32'b00111111011000010101100101110011;
end
if( x >= 32'b01000000000000000000000000000000 && x < 32'b01000000000000001010001111010111)
begin
	y_temp <= 32'b00111111011000011001111001000010;
end
if( x >= 32'b01000000000000001010001111010111 && x < 32'b01000000000000010100011110101110)
begin
	y_temp <= 32'b00111111011000011110001010001011;
end
if( x >= 32'b01000000000000010100011110101110 && x < 32'b01000000000000011110101110000101)
begin
	y_temp <= 32'b00111111011000100010011001001111;
end
if( x >= 32'b01000000000000011110101110000101 && x < 32'b01000000000000101000111101011100)
begin
	y_temp <= 32'b00111111011000100110100110001110;
end
if( x >= 32'b01000000000000101000111101011100 && x < 32'b01000000000000110011001100110011)
begin
	y_temp <= 32'b00111111011000101010110001001010;
end
if( x >= 32'b01000000000000110011001100110011 && x < 32'b01000000000000111101011100001010)
begin
	y_temp <= 32'b00111111011000101110111010000010;
end
if( x >= 32'b01000000000000111101011100001010 && x < 32'b01000000000001000111101011100001)
begin
	y_temp <= 32'b00111111011000110011000000111000;
end
if( x >= 32'b01000000000001000111101011100001 && x < 32'b01000000000001010001111010111000)
begin
	y_temp <= 32'b00111111011000110111000101101100;
end
if( x >= 32'b01000000000001010001111010111000 && x < 32'b01000000000001011100001010001111)
begin
	y_temp <= 32'b00111111011000111011001000011111;
end
if( x >= 32'b01000000000001011100001010001111 && x < 32'b01000000000001100110011001100110)
begin
	y_temp <= 32'b00111111011000111111001001010010;
end
if( x >= 32'b01000000000001100110011001100110 && x < 32'b01000000000001110000101000111101)
begin
	y_temp <= 32'b00111111011001000011001000000100;
end
if( x >= 32'b01000000000001110000101000111101 && x < 32'b01000000000001111010111000010100)
begin
	y_temp <= 32'b00111111011001000111000100111000;
end
if( x >= 32'b01000000000001111010111000010100 && x < 32'b01000000000010000101000111101100)
begin
	y_temp <= 32'b00111111011001001010111111101101;
end
if( x >= 32'b01000000000010000101000111101100 && x < 32'b01000000000010001111010111000011)
begin
	y_temp <= 32'b00111111011001001110111000100100;
end
if( x >= 32'b01000000000010001111010111000011 && x < 32'b01000000000010011001100110011010)
begin
	y_temp <= 32'b00111111011001010010101111011110;
end
if( x >= 32'b01000000000010011001100110011010 && x < 32'b01000000000010100011110101110001)
begin
	y_temp <= 32'b00111111011001010110100100011100;
end
if( x >= 32'b01000000000010100011110101110001 && x < 32'b01000000000010101110000101001000)
begin
	y_temp <= 32'b00111111011001011010010111011110;
end
if( x >= 32'b01000000000010101110000101001000 && x < 32'b01000000000010111000010100011111)
begin
	y_temp <= 32'b00111111011001011110001000100101;
end
if( x >= 32'b01000000000010111000010100011111 && x < 32'b01000000000011000010100011110110)
begin
	y_temp <= 32'b00111111011001100001110111110001;
end
if( x >= 32'b01000000000011000010100011110110 && x < 32'b01000000000011001100110011001101)
begin
	y_temp <= 32'b00111111011001100101100101000100;
end
if( x >= 32'b01000000000011001100110011001101 && x < 32'b01000000000011010111000010100100)
begin
	y_temp <= 32'b00111111011001101001010000011110;
end
if( x >= 32'b01000000000011010111000010100100 && x < 32'b01000000000011100001010001111011)
begin
	y_temp <= 32'b00111111011001101100111010000000;
end
if( x >= 32'b01000000000011100001010001111011 && x < 32'b01000000000011101011100001010010)
begin
	y_temp <= 32'b00111111011001110000100001101010;
end
if( x >= 32'b01000000000011101011100001010010 && x < 32'b01000000000011110101110000101001)
begin
	y_temp <= 32'b00111111011001110100000111011110;
end
if( x >= 32'b01000000000011110101110000101001 && x < 32'b01000000000100000000000000000000)
begin
	y_temp <= 32'b00111111011001110111101011011011;
end
if( x >= 32'b01000000000100000000000000000000 && x < 32'b01000000000100001010001111010111)
begin
	y_temp <= 32'b00111111011001111011001101100011;
end
if( x >= 32'b01000000000100001010001111010111 && x < 32'b01000000000100010100011110101110)
begin
	y_temp <= 32'b00111111011001111110101101110110;
end
if( x >= 32'b01000000000100010100011110101110 && x < 32'b01000000000100011110101110000101)
begin
	y_temp <= 32'b00111111011010000010001100010100;
end
if( x >= 32'b01000000000100011110101110000101 && x < 32'b01000000000100101000111101011100)
begin
	y_temp <= 32'b00111111011010000101101001000000;
end
if( x >= 32'b01000000000100101000111101011100 && x < 32'b01000000000100110011001100110011)
begin
	y_temp <= 32'b00111111011010001001000011111001;
end
if( x >= 32'b01000000000100110011001100110011 && x < 32'b01000000000100111101011100001010)
begin
	y_temp <= 32'b00111111011010001100011101000000;
end
if( x >= 32'b01000000000100111101011100001010 && x < 32'b01000000000101000111101011100001)
begin
	y_temp <= 32'b00111111011010001111110100010101;
end
if( x >= 32'b01000000000101000111101011100001 && x < 32'b01000000000101010001111010111000)
begin
	y_temp <= 32'b00111111011010010011001001111010;
end
if( x >= 32'b01000000000101010001111010111000 && x < 32'b01000000000101011100001010001111)
begin
	y_temp <= 32'b00111111011010010110011101101111;
end
if( x >= 32'b01000000000101011100001010001111 && x < 32'b01000000000101100110011001100110)
begin
	y_temp <= 32'b00111111011010011001101111110101;
end
if( x >= 32'b01000000000101100110011001100110 && x < 32'b01000000000101110000101000111101)
begin
	y_temp <= 32'b00111111011010011101000000001101;
end
if( x >= 32'b01000000000101110000101000111101 && x < 32'b01000000000101111010111000010100)
begin
	y_temp <= 32'b00111111011010100000001110110110;
end
if( x >= 32'b01000000000101111010111000010100 && x < 32'b01000000000110000101000111101100)
begin
	y_temp <= 32'b00111111011010100011011011110011;
end
if( x >= 32'b01000000000110000101000111101100 && x < 32'b01000000000110001111010111000011)
begin
	y_temp <= 32'b00111111011010100110100111000011;
end
if( x >= 32'b01000000000110001111010111000011 && x < 32'b01000000000110011001100110011010)
begin
	y_temp <= 32'b00111111011010101001110000101000;
end
if( x >= 32'b01000000000110011001100110011010 && x < 32'b01000000000110100011110101110001)
begin
	y_temp <= 32'b00111111011010101100111000100001;
end
if( x >= 32'b01000000000110100011110101110001 && x < 32'b01000000000110101110000101001000)
begin
	y_temp <= 32'b00111111011010101111111110110000;
end
if( x >= 32'b01000000000110101110000101001000 && x < 32'b01000000000110111000010100011111)
begin
	y_temp <= 32'b00111111011010110011000011010110;
end
if( x >= 32'b01000000000110111000010100011111 && x < 32'b01000000000111000010100011110110)
begin
	y_temp <= 32'b00111111011010110110000110010011;
end
if( x >= 32'b01000000000111000010100011110110 && x < 32'b01000000000111001100110011001101)
begin
	y_temp <= 32'b00111111011010111001000111100111;
end
if( x >= 32'b01000000000111001100110011001101 && x < 32'b01000000000111010111000010100100)
begin
	y_temp <= 32'b00111111011010111100000111010100;
end
if( x >= 32'b01000000000111010111000010100100 && x < 32'b01000000000111100001010001111011)
begin
	y_temp <= 32'b00111111011010111111000101011010;
end
if( x >= 32'b01000000000111100001010001111011 && x < 32'b01000000000111101011100001010010)
begin
	y_temp <= 32'b00111111011011000010000001111010;
end
if( x >= 32'b01000000000111101011100001010010 && x < 32'b01000000000111110101110000101001)
begin
	y_temp <= 32'b00111111011011000100111100110100;
end
if( x >= 32'b01000000000111110101110000101001 && x < 32'b01000000001000000000000000000000)
begin
	y_temp <= 32'b00111111011011000111110110001010;
end
if( x >= 32'b01000000001000000000000000000000 && x < 32'b01000000001000001010001111010111)
begin
	y_temp <= 32'b00111111011011001010101101111011;
end
if( x >= 32'b01000000001000001010001111010111 && x < 32'b01000000001000010100011110101110)
begin
	y_temp <= 32'b00111111011011001101100100001001;
end
if( x >= 32'b01000000001000010100011110101110 && x < 32'b01000000001000011110101110000101)
begin
	y_temp <= 32'b00111111011011010000011000110101;
end
if( x >= 32'b01000000001000011110101110000101 && x < 32'b01000000001000101000111101011100)
begin
	y_temp <= 32'b00111111011011010011001011111110;
end
if( x >= 32'b01000000001000101000111101011100 && x < 32'b01000000001000110011001100110011)
begin
	y_temp <= 32'b00111111011011010101111101100110;
end
if( x >= 32'b01000000001000110011001100110011 && x < 32'b01000000001000111101011100001010)
begin
	y_temp <= 32'b00111111011011011000101101101101;
end
if( x >= 32'b01000000001000111101011100001010 && x < 32'b01000000001001000111101011100001)
begin
	y_temp <= 32'b00111111011011011011011100010100;
end
if( x >= 32'b01000000001001000111101011100001 && x < 32'b01000000001001010001111010111000)
begin
	y_temp <= 32'b00111111011011011110001001011011;
end
if( x >= 32'b01000000001001010001111010111000 && x < 32'b01000000001001011100001010001111)
begin
	y_temp <= 32'b00111111011011100000110101000100;
end
if( x >= 32'b01000000001001011100001010001111 && x < 32'b01000000001001100110011001100110)
begin
	y_temp <= 32'b00111111011011100011011111001111;
end
if( x >= 32'b01000000001001100110011001100110 && x < 32'b01000000001001110000101000111101)
begin
	y_temp <= 32'b00111111011011100110000111111101;
end
if( x >= 32'b01000000001001110000101000111101 && x < 32'b01000000001001111010111000010100)
begin
	y_temp <= 32'b00111111011011101000101111001110;
end
if( x >= 32'b01000000001001111010111000010100 && x < 32'b01000000001010000101000111101100)
begin
	y_temp <= 32'b00111111011011101011010101000011;
end
if( x >= 32'b01000000001010000101000111101100 && x < 32'b01000000001010001111010111000011)
begin
	y_temp <= 32'b00111111011011101101111001011100;
end
if( x >= 32'b01000000001010001111010111000011 && x < 32'b01000000001010011001100110011010)
begin
	y_temp <= 32'b00111111011011110000011100011011;
end
if( x >= 32'b01000000001010011001100110011010 && x < 32'b01000000001010100011110101110001)
begin
	y_temp <= 32'b00111111011011110010111101111111;
end
if( x >= 32'b01000000001010100011110101110001 && x < 32'b01000000001010101110000101001000)
begin
	y_temp <= 32'b00111111011011110101011110001010;
end
if( x >= 32'b01000000001010101110000101001000 && x < 32'b01000000001010111000010100011111)
begin
	y_temp <= 32'b00111111011011110111111100111101;
end
if( x >= 32'b01000000001010111000010100011111 && x < 32'b01000000001011000010100011110110)
begin
	y_temp <= 32'b00111111011011111010011010010111;
end
if( x >= 32'b01000000001011000010100011110110 && x < 32'b01000000001011001100110011001101)
begin
	y_temp <= 32'b00111111011011111100110110011010;
end
if( x >= 32'b01000000001011001100110011001101 && x < 32'b01000000001011010111000010100100)
begin
	y_temp <= 32'b00111111011011111111010001000110;
end
if( x >= 32'b01000000001011010111000010100100 && x < 32'b01000000001011100001010001111011)
begin
	y_temp <= 32'b00111111011100000001101010011011;
end
if( x >= 32'b01000000001011100001010001111011 && x < 32'b01000000001011101011100001010010)
begin
	y_temp <= 32'b00111111011100000100000010011011;
end
if( x >= 32'b01000000001011101011100001010010 && x < 32'b01000000001011110101110000101001)
begin
	y_temp <= 32'b00111111011100000110011001000110;
end
if( x >= 32'b01000000001011110101110000101001 && x < 32'b01000000001100000000000000000000)
begin
	y_temp <= 32'b00111111011100001000101110011101;
end
if( x >= 32'b01000000001100000000000000000000 && x < 32'b01000000001100001010001111010111)
begin
	y_temp <= 32'b00111111011100001011000010100000;
end
if( x >= 32'b01000000001100001010001111010111 && x < 32'b01000000001100010100011110101110)
begin
	y_temp <= 32'b00111111011100001101010101010001;
end
if( x >= 32'b01000000001100010100011110101110 && x < 32'b01000000001100011110101110000101)
begin
	y_temp <= 32'b00111111011100001111100110101110;
end
if( x >= 32'b01000000001100011110101110000101 && x < 32'b01000000001100101000111101011100)
begin
	y_temp <= 32'b00111111011100010001110110111010;
end
if( x >= 32'b01000000001100101000111101011100 && x < 32'b01000000001100110011001100110011)
begin
	y_temp <= 32'b00111111011100010100000101110101;
end
if( x >= 32'b01000000001100110011001100110011 && x < 32'b01000000001100111101011100001010)
begin
	y_temp <= 32'b00111111011100010110010011011111;
end
if( x >= 32'b01000000001100111101011100001010 && x < 32'b01000000001101000111101011100001)
begin
	y_temp <= 32'b00111111011100011000011111111001;
end
if( x >= 32'b01000000001101000111101011100001 && x < 32'b01000000001101010001111010111000)
begin
	y_temp <= 32'b00111111011100011010101011000100;
end
if( x >= 32'b01000000001101010001111010111000 && x < 32'b01000000001101011100001010001111)
begin
	y_temp <= 32'b00111111011100011100110101000000;
end
if( x >= 32'b01000000001101011100001010001111 && x < 32'b01000000001101100110011001100110)
begin
	y_temp <= 32'b00111111011100011110111101101110;
end
if( x >= 32'b01000000001101100110011001100110 && x < 32'b01000000001101110000101000111101)
begin
	y_temp <= 32'b00111111011100100001000101001110;
end
if( x >= 32'b01000000001101110000101000111101 && x < 32'b01000000001101111010111000010100)
begin
	y_temp <= 32'b00111111011100100011001011100010;
end
if( x >= 32'b01000000001101111010111000010100 && x < 32'b01000000001110000101000111101100)
begin
	y_temp <= 32'b00111111011100100101010000101001;
end
if( x >= 32'b01000000001110000101000111101100 && x < 32'b01000000001110001111010111000011)
begin
	y_temp <= 32'b00111111011100100111010100100100;
end
if( x >= 32'b01000000001110001111010111000011 && x < 32'b01000000001110011001100110011010)
begin
	y_temp <= 32'b00111111011100101001010111010100;
end
if( x >= 32'b01000000001110011001100110011010 && x < 32'b01000000001110100011110101110001)
begin
	y_temp <= 32'b00111111011100101011011000111010;
end
if( x >= 32'b01000000001110100011110101110001 && x < 32'b01000000001110101110000101001000)
begin
	y_temp <= 32'b00111111011100101101011001010110;
end
if( x >= 32'b01000000001110101110000101001000 && x < 32'b01000000001110111000010100011111)
begin
	y_temp <= 32'b00111111011100101111011000101000;
end
if( x >= 32'b01000000001110111000010100011111 && x < 32'b01000000001111000010100011110110)
begin
	y_temp <= 32'b00111111011100110001010110110001;
end
if( x >= 32'b01000000001111000010100011110110 && x < 32'b01000000001111001100110011001101)
begin
	y_temp <= 32'b00111111011100110011010011110010;
end
if( x >= 32'b01000000001111001100110011001101 && x < 32'b01000000001111010111000010100100)
begin
	y_temp <= 32'b00111111011100110101001111101100;
end
if( x >= 32'b01000000001111010111000010100100 && x < 32'b01000000001111100001010001111011)
begin
	y_temp <= 32'b00111111011100110111001010011110;
end
if( x >= 32'b01000000001111100001010001111011 && x < 32'b01000000001111101011100001010010)
begin
	y_temp <= 32'b00111111011100111001000100001010;
end
if( x >= 32'b01000000001111101011100001010010 && x < 32'b01000000001111110101110000101001)
begin
	y_temp <= 32'b00111111011100111010111100101111;
end
if( x >= 32'b01000000001111110101110000101001 && x < 32'b01000000010000000000000000000000)
begin
	y_temp <= 32'b00111111011100111100110100010000;
end
if( x >= 32'b01000000010000000000000000000000 && x < 32'b01000000010000001010001111010111)
begin
	y_temp <= 32'b00111111011100111110101010101011;
end
if( x >= 32'b01000000010000001010001111010111 && x < 32'b01000000010000010100011110101110)
begin
	y_temp <= 32'b00111111011101000000100000000010;
end
if( x >= 32'b01000000010000010100011110101110 && x < 32'b01000000010000011110101110000101)
begin
	y_temp <= 32'b00111111011101000010010100010101;
end
if( x >= 32'b01000000010000011110101110000101 && x < 32'b01000000010000101000111101011100)
begin
	y_temp <= 32'b00111111011101000100000111100101;
end
if( x >= 32'b01000000010000101000111101011100 && x < 32'b01000000010000110011001100110011)
begin
	y_temp <= 32'b00111111011101000101111001110011;
end
if( x >= 32'b01000000010000110011001100110011 && x < 32'b01000000010000111101011100001010)
begin
	y_temp <= 32'b00111111011101000111101010111110;
end
if( x >= 32'b01000000010000111101011100001010 && x < 32'b01000000010001000111101011100001)
begin
	y_temp <= 32'b00111111011101001001011011001000;
end
if( x >= 32'b01000000010001000111101011100001 && x < 32'b01000000010001010001111010111000)
begin
	y_temp <= 32'b00111111011101001011001010010000;
end
if( x >= 32'b01000000010001010001111010111000 && x < 32'b01000000010001011100001010001111)
begin
	y_temp <= 32'b00111111011101001100111000011000;
end
if( x >= 32'b01000000010001011100001010001111 && x < 32'b01000000010001100110011001100110)
begin
	y_temp <= 32'b00111111011101001110100101100000;
end
if( x >= 32'b01000000010001100110011001100110 && x < 32'b01000000010001110000101000111101)
begin
	y_temp <= 32'b00111111011101010000010001101001;
end
if( x >= 32'b01000000010001110000101000111101 && x < 32'b01000000010001111010111000010100)
begin
	y_temp <= 32'b00111111011101010001111100110010;
end
if( x >= 32'b01000000010001111010111000010100 && x < 32'b01000000010010000101000111101100)
begin
	y_temp <= 32'b00111111011101010011100110111101;
end
if( x >= 32'b01000000010010000101000111101100 && x < 32'b01000000010010001111010111000011)
begin
	y_temp <= 32'b00111111011101010101010000001010;
end
if( x >= 32'b01000000010010001111010111000011 && x < 32'b01000000010010011001100110011010)
begin
	y_temp <= 32'b00111111011101010110111000011010;
end
if( x >= 32'b01000000010010011001100110011010 && x < 32'b01000000010010100011110101110001)
begin
	y_temp <= 32'b00111111011101011000011111101101;
end
if( x >= 32'b01000000010010100011110101110001 && x < 32'b01000000010010101110000101001000)
begin
	y_temp <= 32'b00111111011101011010000110000011;
end
if( x >= 32'b01000000010010101110000101001000 && x < 32'b01000000010010111000010100011111)
begin
	y_temp <= 32'b00111111011101011011101011011101;
end
if( x >= 32'b01000000010010111000010100011111 && x < 32'b01000000010011000010100011110110)
begin
	y_temp <= 32'b00111111011101011101001111111100;
end
if( x >= 32'b01000000010011000010100011110110 && x < 32'b01000000010011001100110011001101)
begin
	y_temp <= 32'b00111111011101011110110011100000;
end
if( x >= 32'b01000000010011001100110011001101 && x < 32'b01000000010011010111000010100100)
begin
	y_temp <= 32'b00111111011101100000010110001010;
end
if( x >= 32'b01000000010011010111000010100100 && x < 32'b01000000010011100001010001111011)
begin
	y_temp <= 32'b00111111011101100001110111111001;
end
if( x >= 32'b01000000010011100001010001111011 && x < 32'b01000000010011101011100001010010)
begin
	y_temp <= 32'b00111111011101100011011000110000;
end
if( x >= 32'b01000000010011101011100001010010 && x < 32'b01000000010011110101110000101001)
begin
	y_temp <= 32'b00111111011101100100111000101101;
end
if( x >= 32'b01000000010011110101110000101001 && x < 32'b01000000010100000000000000000000)
begin
	y_temp <= 32'b00111111011101100110010111110001;
end
if( x >= 32'b01000000010100000000000000000000 && x < 32'b01000000010100001010001111010111)
begin
	y_temp <= 32'b00111111011101100111110101111110;
end
if( x >= 32'b01000000010100001010001111010111 && x < 32'b01000000010100010100011110101110)
begin
	y_temp <= 32'b00111111011101101001010011010011;
end
if( x >= 32'b01000000010100010100011110101110 && x < 32'b01000000010100011110101110000101)
begin
	y_temp <= 32'b00111111011101101010101111110001;
end
if( x >= 32'b01000000010100011110101110000101 && x < 32'b01000000010100101000111101011100)
begin
	y_temp <= 32'b00111111011101101100001011011001;
end
if( x >= 32'b01000000010100101000111101011100 && x < 32'b01000000010100110011001100110011)
begin
	y_temp <= 32'b00111111011101101101100110001010;
end
if( x >= 32'b01000000010100110011001100110011 && x < 32'b01000000010100111101011100001010)
begin
	y_temp <= 32'b00111111011101101111000000000110;
end
if( x >= 32'b01000000010100111101011100001010 && x < 32'b01000000010101000111101011100001)
begin
	y_temp <= 32'b00111111011101110000011001001100;
end
if( x >= 32'b01000000010101000111101011100001 && x < 32'b01000000010101010001111010111000)
begin
	y_temp <= 32'b00111111011101110001110001011110;
end
if( x >= 32'b01000000010101010001111010111000 && x < 32'b01000000010101011100001010001111)
begin
	y_temp <= 32'b00111111011101110011001000111011;
end
if( x >= 32'b01000000010101011100001010001111 && x < 32'b01000000010101100110011001100110)
begin
	y_temp <= 32'b00111111011101110100011111100100;
end
if( x >= 32'b01000000010101100110011001100110 && x < 32'b01000000010101110000101000111101)
begin
	y_temp <= 32'b00111111011101110101110101011010;
end
if( x >= 32'b01000000010101110000101000111101 && x < 32'b01000000010101111010111000010100)
begin
	y_temp <= 32'b00111111011101110111001010011101;
end
if( x >= 32'b01000000010101111010111000010100 && x < 32'b01000000010110000101000111101100)
begin
	y_temp <= 32'b00111111011101111000011110101101;
end
if( x >= 32'b01000000010110000101000111101100 && x < 32'b01000000010110001111010111000011)
begin
	y_temp <= 32'b00111111011101111001110010001100;
end
if( x >= 32'b01000000010110001111010111000011 && x < 32'b01000000010110011001100110011010)
begin
	y_temp <= 32'b00111111011101111011000100111000;
end
if( x >= 32'b01000000010110011001100110011010 && x < 32'b01000000010110100011110101110001)
begin
	y_temp <= 32'b00111111011101111100010110110100;
end
if( x >= 32'b01000000010110100011110101110001 && x < 32'b01000000010110101110000101001000)
begin
	y_temp <= 32'b00111111011101111101100111111110;
end
if( x >= 32'b01000000010110101110000101001000 && x < 32'b01000000010110111000010100011111)
begin
	y_temp <= 32'b00111111011101111110111000011000;
end
if( x >= 32'b01000000010110111000010100011111 && x < 32'b01000000010111000010100011110110)
begin
	y_temp <= 32'b00111111011110000000001000000010;
end
if( x >= 32'b01000000010111000010100011110110 && x < 32'b01000000010111001100110011001101)
begin
	y_temp <= 32'b00111111011110000001010110111101;
end
if( x >= 32'b01000000010111001100110011001101 && x < 32'b01000000010111010111000010100100)
begin
	y_temp <= 32'b00111111011110000010100101001000;
end
if( x >= 32'b01000000010111010111000010100100 && x < 32'b01000000010111100001010001111011)
begin
	y_temp <= 32'b00111111011110000011110010100101;
end
if( x >= 32'b01000000010111100001010001111011 && x < 32'b01000000010111101011100001010010)
begin
	y_temp <= 32'b00111111011110000100111111010011;
end
if( x >= 32'b01000000010111101011100001010010 && x < 32'b01000000010111110101110000101001)
begin
	y_temp <= 32'b00111111011110000110001011010011;
end
if( x >= 32'b01000000010111110101110000101001 && x < 32'b01000000011000000000000000000000)
begin
	y_temp <= 32'b00111111011110000111010110100110;
end
if( x >= 32'b01000000011000000000000000000000 && x < 32'b01000000011000001010001111010111)
begin
	y_temp <= 32'b00111111011110001000100001001100;
end
if( x >= 32'b01000000011000001010001111010111 && x < 32'b01000000011000010100011110101110)
begin
	y_temp <= 32'b00111111011110001001101011000100;
end
if( x >= 32'b01000000011000010100011110101110 && x < 32'b01000000011000011110101110000101)
begin
	y_temp <= 32'b00111111011110001010110100010001;
end
if( x >= 32'b01000000011000011110101110000101 && x < 32'b01000000011000101000111101011100)
begin
	y_temp <= 32'b00111111011110001011111100110010;
end
if( x >= 32'b01000000011000101000111101011100 && x < 32'b01000000011000110011001100110011)
begin
	y_temp <= 32'b00111111011110001101000100100111;
end
if( x >= 32'b01000000011000110011001100110011 && x < 32'b01000000011000111101011100001010)
begin
	y_temp <= 32'b00111111011110001110001011110000;
end
if( x >= 32'b01000000011000111101011100001010 && x < 32'b01000000011001000111101011100001)
begin
	y_temp <= 32'b00111111011110001111010010010000;
end
if( x >= 32'b01000000011001000111101011100001 && x < 32'b01000000011001010001111010111000)
begin
	y_temp <= 32'b00111111011110010000011000000100;
end
if( x >= 32'b01000000011001010001111010111000 && x < 32'b01000000011001011100001010001111)
begin
	y_temp <= 32'b00111111011110010001011101001111;
end
if( x >= 32'b01000000011001011100001010001111 && x < 32'b01000000011001100110011001100110)
begin
	y_temp <= 32'b00111111011110010010100001110000;
end
if( x >= 32'b01000000011001100110011001100110 && x < 32'b01000000011001110000101000111101)
begin
	y_temp <= 32'b00111111011110010011100101100111;
end
if( x >= 32'b01000000011001110000101000111101 && x < 32'b01000000011001111010111000010100)
begin
	y_temp <= 32'b00111111011110010100101000110110;
end
if( x >= 32'b01000000011001111010111000010100 && x < 32'b01000000011010000101000111101100)
begin
	y_temp <= 32'b00111111011110010101101011011100;
end
if( x >= 32'b01000000011010000101000111101100 && x < 32'b01000000011010001111010111000011)
begin
	y_temp <= 32'b00111111011110010110101101011010;
end
if( x >= 32'b01000000011010001111010111000011 && x < 32'b01000000011010011001100110011010)
begin
	y_temp <= 32'b00111111011110010111101110110000;
end
if( x >= 32'b01000000011010011001100110011010 && x < 32'b01000000011010100011110101110001)
begin
	y_temp <= 32'b00111111011110011000101111011110;
end
if( x >= 32'b01000000011010100011110101110001 && x < 32'b01000000011010101110000101001000)
begin
	y_temp <= 32'b00111111011110011001101111100101;
end
if( x >= 32'b01000000011010101110000101001000 && x < 32'b01000000011010111000010100011111)
begin
	y_temp <= 32'b00111111011110011010101111000110;
end
if( x >= 32'b01000000011010111000010100011111 && x < 32'b01000000011011000010100011110110)
begin
	y_temp <= 32'b00111111011110011011101110000000;
end
if( x >= 32'b01000000011011000010100011110110 && x < 32'b01000000011011001100110011001101)
begin
	y_temp <= 32'b00111111011110011100101100010100;
end
if( x >= 32'b01000000011011001100110011001101 && x < 32'b01000000011011010111000010100100)
begin
	y_temp <= 32'b00111111011110011101101010000010;
end
if( x >= 32'b01000000011011010111000010100100 && x < 32'b01000000011011100001010001111011)
begin
	y_temp <= 32'b00111111011110011110100111001011;
end
if( x >= 32'b01000000011011100001010001111011 && x < 32'b01000000011011101011100001010010)
begin
	y_temp <= 32'b00111111011110011111100011101111;
end
if( x >= 32'b01000000011011101011100001010010 && x < 32'b01000000011011110101110000101001)
begin
	y_temp <= 32'b00111111011110100000011111101110;
end
if( x >= 32'b01000000011011110101110000101001 && x < 32'b01000000011100000000000000000000)
begin
	y_temp <= 32'b00111111011110100001011011001000;
end
if( x >= 32'b01000000011100000000000000000000 && x < 32'b01000000011100001010001111010111)
begin
	y_temp <= 32'b00111111011110100010010101111110;
end
if( x >= 32'b01000000011100001010001111010111 && x < 32'b01000000011100010100011110101110)
begin
	y_temp <= 32'b00111111011110100011010000010001;
end
if( x >= 32'b01000000011100010100011110101110 && x < 32'b01000000011100011110101110000101)
begin
	y_temp <= 32'b00111111011110100100001010000000;
end
if( x >= 32'b01000000011100011110101110000101 && x < 32'b01000000011100101000111101011100)
begin
	y_temp <= 32'b00111111011110100101000011001100;
end
if( x >= 32'b01000000011100101000111101011100 && x < 32'b01000000011100110011001100110011)
begin
	y_temp <= 32'b00111111011110100101111011110110;
end
if( x >= 32'b01000000011100110011001100110011 && x < 32'b01000000011100111101011100001010)
begin
	y_temp <= 32'b00111111011110100110110011111100;
end
if( x >= 32'b01000000011100111101011100001010 && x < 32'b01000000011101000111101011100001)
begin
	y_temp <= 32'b00111111011110100111101011100001;
end
if( x >= 32'b01000000011101000111101011100001 && x < 32'b01000000011101010001111010111000)
begin
	y_temp <= 32'b00111111011110101000100010100100;
end
if( x >= 32'b01000000011101010001111010111000 && x < 32'b01000000011101011100001010001111)
begin
	y_temp <= 32'b00111111011110101001011001000101;
end
if( x >= 32'b01000000011101011100001010001111 && x < 32'b01000000011101100110011001100110)
begin
	y_temp <= 32'b00111111011110101010001111000101;
end
if( x >= 32'b01000000011101100110011001100110 && x < 32'b01000000011101110000101000111101)
begin
	y_temp <= 32'b00111111011110101011000100100100;
end
if( x >= 32'b01000000011101110000101000111101 && x < 32'b01000000011101111010111000010100)
begin
	y_temp <= 32'b00111111011110101011111001100010;
end
if( x >= 32'b01000000011101111010111000010100 && x < 32'b01000000011110000101000111101100)
begin
	y_temp <= 32'b00111111011110101100101110000000;
end
if( x >= 32'b01000000011110000101000111101100 && x < 32'b01000000011110001111010111000011)
begin
	y_temp <= 32'b00111111011110101101100001111110;
end
if( x >= 32'b01000000011110001111010111000011 && x < 32'b01000000011110011001100110011010)
begin
	y_temp <= 32'b00111111011110101110010101011100;
end
if( x >= 32'b01000000011110011001100110011010 && x < 32'b01000000011110100011110101110001)
begin
	y_temp <= 32'b00111111011110101111001000011010;
end
if( x >= 32'b01000000011110100011110101110001 && x < 32'b01000000011110101110000101001000)
begin
	y_temp <= 32'b00111111011110101111111010111010;
end
if( x >= 32'b01000000011110101110000101001000 && x < 32'b01000000011110111000010100011111)
begin
	y_temp <= 32'b00111111011110110000101100111010;
end
if( x >= 32'b01000000011110111000010100011111 && x < 32'b01000000011111000010100011110110)
begin
	y_temp <= 32'b00111111011110110001011110011100;
end
if( x >= 32'b01000000011111000010100011110110 && x < 32'b01000000011111001100110011001101)
begin
	y_temp <= 32'b00111111011110110010001111100000;
end
if( x >= 32'b01000000011111001100110011001101 && x < 32'b01000000011111010111000010100100)
begin
	y_temp <= 32'b00111111011110110011000000000101;
end
if( x >= 32'b01000000011111010111000010100100 && x < 32'b01000000011111100001010001111011)
begin
	y_temp <= 32'b00111111011110110011110000001101;
end
if( x >= 32'b01000000011111100001010001111011 && x < 32'b01000000011111101011100001010010)
begin
	y_temp <= 32'b00111111011110110100011111110111;
end
if( x >= 32'b01000000011111101011100001010010 && x < 32'b01000000011111110101110000101001)
begin
	y_temp <= 32'b00111111011110110101001111000100;
end
if( x >= 32'b01000000011111110101110000101001 && x < 32'b01000000100000000000000000000000)
begin
	y_temp <= 32'b00111111011110110101111101110100;
end
if( x >= 32'b01000000100000000000000000000000 && x < 32'b01000000100000000101000111101100)
begin
	y_temp <= 32'b00111111011110110110101100001000;
end
if( x >= 32'b01000000100000000101000111101100 && x < 32'b01000000100000001010001111010111)
begin
	y_temp <= 32'b00111111011110110111011001111110;
end
if( x >= 32'b01000000100000001010001111010111 && x < 32'b01000000100000001111010111000011)
begin
	y_temp <= 32'b00111111011110111000000111011001;
end
if( x >= 32'b01000000100000001111010111000011 && x < 32'b01000000100000010100011110101110)
begin
	y_temp <= 32'b00111111011110111000110100011000;
end
if( x >= 32'b01000000100000010100011110101110 && x < 32'b01000000100000011001100110011010)
begin
	y_temp <= 32'b00111111011110111001100000111011;
end
if( x >= 32'b01000000100000011001100110011010 && x < 32'b01000000100000011110101110000101)
begin
	y_temp <= 32'b00111111011110111010001101000011;
end
if( x >= 32'b01000000100000011110101110000101 && x < 32'b01000000100000100011110101110001)
begin
	y_temp <= 32'b00111111011110111010111000101111;
end
if( x >= 32'b01000000100000100011110101110001 && x < 32'b01000000100000101000111101011100)
begin
	y_temp <= 32'b00111111011110111011100100000001;
end
if( x >= 32'b01000000100000101000111101011100 && x < 32'b01000000100000101110000101001000)
begin
	y_temp <= 32'b00111111011110111100001110111000;
end
if( x >= 32'b01000000100000101110000101001000 && x < 32'b01000000100000110011001100110011)
begin
	y_temp <= 32'b00111111011110111100111001010101;
end
if( x >= 32'b01000000100000110011001100110011 && x < 32'b01000000100000111000010100011111)
begin
	y_temp <= 32'b00111111011110111101100011010111;
end
if( x >= 32'b01000000100000111000010100011111 && x < 32'b01000000100000111101011100001010)
begin
	y_temp <= 32'b00111111011110111110001101000000;
end
if( x >= 32'b01000000100000111101011100001010 && x < 32'b01000000100001000010100011110110)
begin
	y_temp <= 32'b00111111011110111110110110001111;
end
if( x >= 32'b01000000100001000010100011110110 && x < 32'b01000000100001000111101011100001)
begin
	y_temp <= 32'b00111111011110111111011111000101;
end
if( x >= 32'b01000000100001000111101011100001 && x < 32'b01000000100001001100110011001101)
begin
	y_temp <= 32'b00111111011111000000000111100001;
end
if( x >= 32'b01000000100001001100110011001101 && x < 32'b01000000100001010001111010111000)
begin
	y_temp <= 32'b00111111011111000000101111100100;
end
if( x >= 32'b01000000100001010001111010111000 && x < 32'b01000000100001010111000010100100)
begin
	y_temp <= 32'b00111111011111000001010111001111;
end
if( x >= 32'b01000000100001010111000010100100 && x < 32'b01000000100001011100001010001111)
begin
	y_temp <= 32'b00111111011111000001111110100001;
end
if( x >= 32'b01000000100001011100001010001111 && x < 32'b01000000100001100001010001111011)
begin
	y_temp <= 32'b00111111011111000010100101011011;
end
if( x >= 32'b01000000100001100001010001111011 && x < 32'b01000000100001100110011001100110)
begin
	y_temp <= 32'b00111111011111000011001011111101;
end
if( x >= 32'b01000000100001100110011001100110 && x < 32'b01000000100001101011100001010010)
begin
	y_temp <= 32'b00111111011111000011110010000111;
end
if( x >= 32'b01000000100001101011100001010010 && x < 32'b01000000100001110000101000111101)
begin
	y_temp <= 32'b00111111011111000100010111111001;
end
if( x >= 32'b01000000100001110000101000111101 && x < 32'b01000000100001110101110000101001)
begin
	y_temp <= 32'b00111111011111000100111101010101;
end
if( x >= 32'b01000000100001110101110000101001 && x < 32'b01000000100001111010111000010100)
begin
	y_temp <= 32'b00111111011111000101100010011000;
end
if( x >= 32'b01000000100001111010111000010100 && x < 32'b01000000100010000000000000000000)
begin
	y_temp <= 32'b00111111011111000110000111000110;
end
if( x >= 32'b01000000100010000000000000000000 && x < 32'b01000000100010000101000111101100)
begin
	y_temp <= 32'b00111111011111000110101011011100;
end
if( x >= 32'b01000000100010000101000111101100 && x < 32'b01000000100010001010001111010111)
begin
	y_temp <= 32'b00111111011111000111001111011100;
end
if( x >= 32'b01000000100010001010001111010111 && x < 32'b01000000100010001111010111000011)
begin
	y_temp <= 32'b00111111011111000111110011000101;
end
if( x >= 32'b01000000100010001111010111000011 && x < 32'b01000000100010010100011110101110)
begin
	y_temp <= 32'b00111111011111001000010110011001;
end
if( x >= 32'b01000000100010010100011110101110 && x < 32'b01000000100010011001100110011010)
begin
	y_temp <= 32'b00111111011111001000111001010110;
end
if( x >= 32'b01000000100010011001100110011010 && x < 32'b01000000100010011110101110000101)
begin
	y_temp <= 32'b00111111011111001001011011111110;
end
if( x >= 32'b01000000100010011110101110000101 && x < 32'b01000000100010100011110101110001)
begin
	y_temp <= 32'b00111111011111001001111110010000;
end
if( x >= 32'b01000000100010100011110101110001 && x < 32'b01000000100010101000111101011100)
begin
	y_temp <= 32'b00111111011111001010100000001110;
end
if( x >= 32'b01000000100010101000111101011100 && x < 32'b01000000100010101110000101001000)
begin
	y_temp <= 32'b00111111011111001011000001110110;
end
if( x >= 32'b01000000100010101110000101001000 && x < 32'b01000000100010110011001100110011)
begin
	y_temp <= 32'b00111111011111001011100011001001;
end
if( x >= 32'b01000000100010110011001100110011 && x < 32'b01000000100010111000010100011111)
begin
	y_temp <= 32'b00111111011111001100000100001000;
end
if( x >= 32'b01000000100010111000010100011111 && x < 32'b01000000100010111101011100001010)
begin
	y_temp <= 32'b00111111011111001100100100110010;
end
if( x >= 32'b01000000100010111101011100001010 && x < 32'b01000000100011000010100011110110)
begin
	y_temp <= 32'b00111111011111001101000101001000;
end
if( x >= 32'b01000000100011000010100011110110 && x < 32'b01000000100011000111101011100001)
begin
	y_temp <= 32'b00111111011111001101100101001001;
end
if( x >= 32'b01000000100011000111101011100001 && x < 32'b01000000100011001100110011001101)
begin
	y_temp <= 32'b00111111011111001110000100110111;
end
if( x >= 32'b01000000100011001100110011001101 && x < 32'b01000000100011010001111010111000)
begin
	y_temp <= 32'b00111111011111001110100100010001;
end
if( x >= 32'b01000000100011010001111010111000 && x < 32'b01000000100011010111000010100100)
begin
	y_temp <= 32'b00111111011111001111000011011000;
end
if( x >= 32'b01000000100011010111000010100100 && x < 32'b01000000100011011100001010001111)
begin
	y_temp <= 32'b00111111011111001111100010001011;
end
if( x >= 32'b01000000100011011100001010001111 && x < 32'b01000000100011100001010001111011)
begin
	y_temp <= 32'b00111111011111010000000000101011;
end
if( x >= 32'b01000000100011100001010001111011 && x < 32'b01000000100011100110011001100110)
begin
	y_temp <= 32'b00111111011111010000011110111000;
end
if( x >= 32'b01000000100011100110011001100110 && x < 32'b01000000100011101011100001010010)
begin
	y_temp <= 32'b00111111011111010000111100110011;
end
if( x >= 32'b01000000100011101011100001010010 && x < 32'b01000000100011110000101000111101)
begin
	y_temp <= 32'b00111111011111010001011010011011;
end
if( x >= 32'b01000000100011110000101000111101 && x < 32'b01000000100011110101110000101001)
begin
	y_temp <= 32'b00111111011111010001110111110000;
end
if( x >= 32'b01000000100011110101110000101001 && x < 32'b01000000100011111010111000010100)
begin
	y_temp <= 32'b00111111011111010010010100110011;
end
if( x >= 32'b01000000100011111010111000010100 && x < 32'b01000000100100000000000000000000)
begin
	y_temp <= 32'b00111111011111010010110001100100;
end
if( x >= 32'b01000000100100000000000000000000 && x < 32'b01000000100100000101000111101100)
begin
	y_temp <= 32'b00111111011111010011001110000011;
end
if( x >= 32'b01000000100100000101000111101100 && x < 32'b01000000100100001010001111010111)
begin
	y_temp <= 32'b00111111011111010011101010010000;
end
if( x >= 32'b01000000100100001010001111010111 && x < 32'b01000000100100001111010111000011)
begin
	y_temp <= 32'b00111111011111010100000110001100;
end
if( x >= 32'b01000000100100001111010111000011 && x < 32'b01000000100100010100011110101110)
begin
	y_temp <= 32'b00111111011111010100100001110110;
end
if( x >= 32'b01000000100100010100011110101110 && x < 32'b01000000100100011001100110011010)
begin
	y_temp <= 32'b00111111011111010100111101001111;
end
if( x >= 32'b01000000100100011001100110011010 && x < 32'b01000000100100011110101110000101)
begin
	y_temp <= 32'b00111111011111010101011000010111;
end
if( x >= 32'b01000000100100011110101110000101 && x < 32'b01000000100100100011110101110001)
begin
	y_temp <= 32'b00111111011111010101110011001111;
end
if( x >= 32'b01000000100100100011110101110001 && x < 32'b01000000100100101000111101011100)
begin
	y_temp <= 32'b00111111011111010110001101110101;
end
if( x >= 32'b01000000100100101000111101011100 && x < 32'b01000000100100101110000101001000)
begin
	y_temp <= 32'b00111111011111010110101000001011;
end
if( x >= 32'b01000000100100101110000101001000 && x < 32'b01000000100100110011001100110011)
begin
	y_temp <= 32'b00111111011111010111000010010000;
end
if( x >= 32'b01000000100100110011001100110011 && x < 32'b01000000100100111000010100011111)
begin
	y_temp <= 32'b00111111011111010111011100000101;
end
if( x >= 32'b01000000100100111000010100011111 && x < 32'b01000000100100111101011100001010)
begin
	y_temp <= 32'b00111111011111010111110101101010;
end
if( x >= 32'b01000000100100111101011100001010 && x < 32'b01000000100101000010100011110110)
begin
	y_temp <= 32'b00111111011111011000001110111111;
end
if( x >= 32'b01000000100101000010100011110110 && x < 32'b01000000100101000111101011100001)
begin
	y_temp <= 32'b00111111011111011000101000000100;
end
if( x >= 32'b01000000100101000111101011100001 && x < 32'b01000000100101001100110011001101)
begin
	y_temp <= 32'b00111111011111011001000000111001;
end
if( x >= 32'b01000000100101001100110011001101 && x < 32'b01000000100101010001111010111000)
begin
	y_temp <= 32'b00111111011111011001011001011111;
end
if( x >= 32'b01000000100101010001111010111000 && x < 32'b01000000100101010111000010100100)
begin
	y_temp <= 32'b00111111011111011001110001110110;
end
if( x >= 32'b01000000100101010111000010100100 && x < 32'b01000000100101011100001010001111)
begin
	y_temp <= 32'b00111111011111011010001001111101;
end
if( x >= 32'b01000000100101011100001010001111 && x < 32'b01000000100101100001010001111011)
begin
	y_temp <= 32'b00111111011111011010100001110101;
end
if( x >= 32'b01000000100101100001010001111011 && x < 32'b01000000100101100110011001100110)
begin
	y_temp <= 32'b00111111011111011010111001011111;
end
if( x >= 32'b01000000100101100110011001100110 && x < 32'b01000000100101101011100001010010)
begin
	y_temp <= 32'b00111111011111011011010000111001;
end
if( x >= 32'b01000000100101101011100001010010 && x < 32'b01000000100101110000101000111101)
begin
	y_temp <= 32'b00111111011111011011101000000101;
end
if( x >= 32'b01000000100101110000101000111101 && x < 32'b01000000100101110101110000101001)
begin
	y_temp <= 32'b00111111011111011011111111000011;
end
if( x >= 32'b01000000100101110101110000101001 && x < 32'b01000000100101111010111000010100)
begin
	y_temp <= 32'b00111111011111011100010101110010;
end
if( x >= 32'b01000000100101111010111000010100 && x < 32'b01000000100110000000000000000000)
begin
	y_temp <= 32'b00111111011111011100101100010011;
end
if( x >= 32'b01000000100110000000000000000000 && x < 32'b01000000100110000101000111101100)
begin
	y_temp <= 32'b00111111011111011101000010100101;
end
if( x >= 32'b01000000100110000101000111101100 && x < 32'b01000000100110001010001111010111)
begin
	y_temp <= 32'b00111111011111011101011000101010;
end
if( x >= 32'b01000000100110001010001111010111 && x < 32'b01000000100110001111010111000011)
begin
	y_temp <= 32'b00111111011111011101101110100001;
end
if( x >= 32'b01000000100110001111010111000011 && x < 32'b01000000100110010100011110101110)
begin
	y_temp <= 32'b00111111011111011110000100001010;
end
if( x >= 32'b01000000100110010100011110101110 && x < 32'b01000000100110011001100110011010)
begin
	y_temp <= 32'b00111111011111011110011001100110;
end
if( x >= 32'b01000000100110011001100110011010 && x < 32'b01000000100110011110101110000101)
begin
	y_temp <= 32'b00111111011111011110101110110100;
end
if( x >= 32'b01000000100110011110101110000101 && x < 32'b01000000100110100011110101110001)
begin
	y_temp <= 32'b00111111011111011111000011110101;
end
if( x >= 32'b01000000100110100011110101110001 && x < 32'b01000000100110101000111101011100)
begin
	y_temp <= 32'b00111111011111011111011000101001;
end
if( x >= 32'b01000000100110101000111101011100 && x < 32'b01000000100110101110000101001000)
begin
	y_temp <= 32'b00111111011111011111101101010000;
end
if( x >= 32'b01000000100110101110000101001000 && x < 32'b01000000100110110011001100110011)
begin
	y_temp <= 32'b00111111011111100000000001101010;
end
if( x >= 32'b01000000100110110011001100110011 && x < 32'b01000000100110111000010100011111)
begin
	y_temp <= 32'b00111111011111100000010101110111;
end
if( x >= 32'b01000000100110111000010100011111 && x < 32'b01000000100110111101011100001010)
begin
	y_temp <= 32'b00111111011111100000101001110111;
end
if( x >= 32'b01000000100110111101011100001010 && x < 32'b01000000100111000010100011110110)
begin
	y_temp <= 32'b00111111011111100000111101101011;
end
if( x >= 32'b01000000100111000010100011110110 && x < 32'b01000000100111000111101011100001)
begin
	y_temp <= 32'b00111111011111100001010001010010;
end
if( x >= 32'b01000000100111000111101011100001 && x < 32'b01000000100111001100110011001101)
begin
	y_temp <= 32'b00111111011111100001100100101110;
end
if( x >= 32'b01000000100111001100110011001101 && x < 32'b01000000100111010001111010111000)
begin
	y_temp <= 32'b00111111011111100001110111111100;
end
if( x >= 32'b01000000100111010001111010111000 && x < 32'b01000000100111010111000010100100)
begin
	y_temp <= 32'b00111111011111100010001010111111;
end
if( x >= 32'b01000000100111010111000010100100 && x < 32'b01000000100111011100001010001111)
begin
	y_temp <= 32'b00111111011111100010011101110110;
end
if( x >= 32'b01000000100111011100001010001111 && x < 32'b01000000100111100001010001111011)
begin
	y_temp <= 32'b00111111011111100010110000100001;
end
if( x >= 32'b01000000100111100001010001111011 && x < 32'b01000000100111100110011001100110)
begin
	y_temp <= 32'b00111111011111100011000011000001;
end
if( x >= 32'b01000000100111100110011001100110 && x < 32'b01000000100111101011100001010010)
begin
	y_temp <= 32'b00111111011111100011010101010100;
end
if( x >= 32'b01000000100111101011100001010010 && x < 32'b01000000100111110000101000111101)
begin
	y_temp <= 32'b00111111011111100011100111011101;
end
if( x >= 32'b01000000100111110000101000111101 && x < 32'b01000000100111110101110000101001)
begin
	y_temp <= 32'b00111111011111100011111001011010;
end
if( x >= 32'b01000000100111110101110000101001 && x < 32'b01000000100111111010111000010100)
begin
	y_temp <= 32'b00111111011111100100001011001011;
end
if( x >= 32'b01000000100111111010111000010100 && x < 32'b01000000101000000000000000000000)
begin
	y_temp <= 32'b00111111011111100100011100110010;
end
if( x >= 32'b01000000101000000000000000000000 )
begin
	y_temp <= 32'b00111111100000000000000000000000;
end
if( x == 0 )
begin
	y_temp <= 32'b00111111000000000000000000000000;
end

end
else
begin
if( x <= 32'b11000000101000000000000000000000 && x > 32'b11000000100111111010111000010100)
begin
	y_temp <= 32'b00111011110111000110011100111011;
end
if( x <= 32'b11000000100111111010111000010100 && x > 32'b11000000100111110101110000101001)
begin
	y_temp <= 32'b00111011110111101001101001110001;
end
if( x <= 32'b11000000100111110101110000101001 && x > 32'b11000000100111110000101000111101)
begin
	y_temp <= 32'b00111011111000001101001100111100;
end
if( x <= 32'b11000000100111110000101000111101 && x > 32'b11000000100111101011100001010010)
begin
	y_temp <= 32'b00111011111000110001000110101011;
end
if( x <= 32'b11000000100111101011100001010010 && x > 32'b11000000100111100110011001100110)
begin
	y_temp <= 32'b00111011111001010101010111001011;
end
if( x <= 32'b11000000100111100110011001100110 && x > 32'b11000000100111100001010001111011)
begin
	y_temp <= 32'b00111011111001111001111110101010;
end
if( x <= 32'b11000000100111100001010001111011 && x > 32'b11000000100111011100001010001111)
begin
	y_temp <= 32'b00111011111010011110111101010111;
end
if( x <= 32'b11000000100111011100001010001111 && x > 32'b11000000100111010111000010100100)
begin
	y_temp <= 32'b00111011111011000100010011100001;
end
if( x <= 32'b11000000100111010111000010100100 && x > 32'b11000000100111010001111010111000)
begin
	y_temp <= 32'b00111011111011101010000001010110;
end
if( x <= 32'b11000000100111010001111010111000 && x > 32'b11000000100111001100110011001101)
begin
	y_temp <= 32'b00111011111100010000000111000100;
end
if( x <= 32'b11000000100111001100110011001101 && x > 32'b11000000100111000111101011100001)
begin
	y_temp <= 32'b00111011111100110110100100111100;
end
if( x <= 32'b11000000100111000111101011100001 && x > 32'b11000000100111000010100011110110)
begin
	y_temp <= 32'b00111011111101011101011011001011;
end
if( x <= 32'b11000000100111000010100011110110 && x > 32'b11000000100110111101011100001010)
begin
	y_temp <= 32'b00111011111110000100101010000010;
end
if( x <= 32'b11000000100110111101011100001010 && x > 32'b11000000100110111000010100011111)
begin
	y_temp <= 32'b00111011111110101100010001101111;
end
if( x <= 32'b11000000100110111000010100011111 && x > 32'b11000000100110110011001100110011)
begin
	y_temp <= 32'b00111011111111010100010010100001;
end
if( x <= 32'b11000000100110110011001100110011 && x > 32'b11000000100110101110000101001000)
begin
	y_temp <= 32'b00111011111111111100101100101010;
end
if( x <= 32'b11000000100110101110000101001000 && x > 32'b11000000100110101000111101011100)
begin
	y_temp <= 32'b00111100000000010010110000001100;
end
if( x <= 32'b11000000100110101000111101011100 && x > 32'b11000000100110100011110101110001)
begin
	y_temp <= 32'b00111100000000100111010110111101;
end
if( x <= 32'b11000000100110100011110101110001 && x > 32'b11000000100110011110101110000101)
begin
	y_temp <= 32'b00111100000000111100001010110001;
end
if( x <= 32'b11000000100110011110101110000101 && x > 32'b11000000100110011001100110011010)
begin
	y_temp <= 32'b00111100000001010001001011110000;
end
if( x <= 32'b11000000100110011001100110011010 && x > 32'b11000000100110010100011110101110)
begin
	y_temp <= 32'b00111100000001100110011010000010;
end
if( x <= 32'b11000000100110010100011110101110 && x > 32'b11000000100110001111010111000011)
begin
	y_temp <= 32'b00111100000001111011110101101111;
end
if( x <= 32'b11000000100110001111010111000011 && x > 32'b11000000100110001010001111010111)
begin
	y_temp <= 32'b00111100000010010001011111000000;
end
if( x <= 32'b11000000100110001010001111010111 && x > 32'b11000000100110000101000111101100)
begin
	y_temp <= 32'b00111100000010100111010101111100;
end
if( x <= 32'b11000000100110000101000111101100 && x > 32'b11000000100110000000000000000000)
begin
	y_temp <= 32'b00111100000010111101011010101110;
end
if( x <= 32'b11000000100110000000000000000000 && x > 32'b11000000100101111010111000010100)
begin
	y_temp <= 32'b00111100000011010011101101011100;
end
if( x <= 32'b11000000100101111010111000010100 && x > 32'b11000000100101110101110000101001)
begin
	y_temp <= 32'b00111100000011101010001110010000;
end
if( x <= 32'b11000000100101110101110000101001 && x > 32'b11000000100101110000101000111101)
begin
	y_temp <= 32'b00111100000100000000111101010011;
end
if( x <= 32'b11000000100101110000101000111101 && x > 32'b11000000100101101011100001010010)
begin
	y_temp <= 32'b00111100000100010111111010101101;
end
if( x <= 32'b11000000100101101011100001010010 && x > 32'b11000000100101100110011001100110)
begin
	y_temp <= 32'b00111100000100101111000110101000;
end
if( x <= 32'b11000000100101100110011001100110 && x > 32'b11000000100101100001010001111011)
begin
	y_temp <= 32'b00111100000101000110100001001011;
end
if( x <= 32'b11000000100101100001010001111011 && x > 32'b11000000100101011100001010001111)
begin
	y_temp <= 32'b00111100000101011110001010100001;
end
if( x <= 32'b11000000100101011100001010001111 && x > 32'b11000000100101010111000010100100)
begin
	y_temp <= 32'b00111100000101110110000010110011;
end
if( x <= 32'b11000000100101010111000010100100 && x > 32'b11000000100101010001111010111000)
begin
	y_temp <= 32'b00111100000110001110001010001001;
end
if( x <= 32'b11000000100101010001111010111000 && x > 32'b11000000100101001100110011001101)
begin
	y_temp <= 32'b00111100000110100110100000101101;
end
if( x <= 32'b11000000100101001100110011001101 && x > 32'b11000000100101000111101011100001)
begin
	y_temp <= 32'b00111100000110111111000110101001;
end
if( x <= 32'b11000000100101000111101011100001 && x > 32'b11000000100101000010100011110110)
begin
	y_temp <= 32'b00111100000111010111111100000110;
end
if( x <= 32'b11000000100101000010100011110110 && x > 32'b11000000100100111101011100001010)
begin
	y_temp <= 32'b00111100000111110001000001001101;
end
if( x <= 32'b11000000100100111101011100001010 && x > 32'b11000000100100111000010100011111)
begin
	y_temp <= 32'b00111100001000001010010110001001;
end
if( x <= 32'b11000000100100111000010100011111 && x > 32'b11000000100100110011001100110011)
begin
	y_temp <= 32'b00111100001000100011111011000011;
end
if( x <= 32'b11000000100100110011001100110011 && x > 32'b11000000100100101110000101001000)
begin
	y_temp <= 32'b00111100001000111101110000000100;
end
if( x <= 32'b11000000100100101110000101001000 && x > 32'b11000000100100101000111101011100)
begin
	y_temp <= 32'b00111100001001010111110101011000;
end
if( x <= 32'b11000000100100101000111101011100 && x > 32'b11000000100100100011110101110001)
begin
	y_temp <= 32'b00111100001001110010001011000111;
end
if( x <= 32'b11000000100100100011110101110001 && x > 32'b11000000100100011110101110000101)
begin
	y_temp <= 32'b00111100001010001100110001011101;
end
if( x <= 32'b11000000100100011110101110000101 && x > 32'b11000000100100011001100110011010)
begin
	y_temp <= 32'b00111100001010100111101000100011;
end
if( x <= 32'b11000000100100011001100110011010 && x > 32'b11000000100100010100011110101110)
begin
	y_temp <= 32'b00111100001011000010110000100011;
end
if( x <= 32'b11000000100100010100011110101110 && x > 32'b11000000100100001111010111000011)
begin
	y_temp <= 32'b00111100001011011110001001101000;
end
if( x <= 32'b11000000100100001111010111000011 && x > 32'b11000000100100001010001111010111)
begin
	y_temp <= 32'b00111100001011111001110011111101;
end
if( x <= 32'b11000000100100001010001111010111 && x > 32'b11000000100100000101000111101100)
begin
	y_temp <= 32'b00111100001100010101101111101101;
end
if( x <= 32'b11000000100100000101000111101100 && x > 32'b11000000100100000000000000000000)
begin
	y_temp <= 32'b00111100001100110001111101000001;
end
if( x <= 32'b11000000100100000000000000000000 && x > 32'b11000000100011111010111000010100)
begin
	y_temp <= 32'b00111100001101001110011100000100;
end
if( x <= 32'b11000000100011111010111000010100 && x > 32'b11000000100011110101110000101001)
begin
	y_temp <= 32'b00111100001101101011001101000011;
end
if( x <= 32'b11000000100011110101110000101001 && x > 32'b11000000100011110000101000111101)
begin
	y_temp <= 32'b00111100001110001000010000000111;
end
if( x <= 32'b11000000100011110000101000111101 && x > 32'b11000000100011101011100001010010)
begin
	y_temp <= 32'b00111100001110100101100101011011;
end
if( x <= 32'b11000000100011101011100001010010 && x > 32'b11000000100011100110011001100110)
begin
	y_temp <= 32'b00111100001111000011001101001100;
end
if( x <= 32'b11000000100011100110011001100110 && x > 32'b11000000100011100001010001111011)
begin
	y_temp <= 32'b00111100001111100001000111100011;
end
if( x <= 32'b11000000100011100001010001111011 && x > 32'b11000000100011011100001010001111)
begin
	y_temp <= 32'b00111100001111111111010100101110;
end
if( x <= 32'b11000000100011011100001010001111 && x > 32'b11000000100011010111000010100100)
begin
	y_temp <= 32'b00111100010000011101110100110110;
end
if( x <= 32'b11000000100011010111000010100100 && x > 32'b11000000100011010001111010111000)
begin
	y_temp <= 32'b00111100010000111100101000001000;
end
if( x <= 32'b11000000100011010001111010111000 && x > 32'b11000000100011001100110011001101)
begin
	y_temp <= 32'b00111100010001011011101110110000;
end
if( x <= 32'b11000000100011001100110011001101 && x > 32'b11000000100011000111101011100001)
begin
	y_temp <= 32'b00111100010001111011001000111001;
end
if( x <= 32'b11000000100011000111101011100001 && x > 32'b11000000100011000010100011110110)
begin
	y_temp <= 32'b00111100010010011010110110110000;
end
if( x <= 32'b11000000100011000010100011110110 && x > 32'b11000000100010111101011100001010)
begin
	y_temp <= 32'b00111100010010111010111000011111;
end
if( x <= 32'b11000000100010111101011100001010 && x > 32'b11000000100010111000010100011111)
begin
	y_temp <= 32'b00111100010011011011001110010101;
end
if( x <= 32'b11000000100010111000010100011111 && x > 32'b11000000100010110011001100110011)
begin
	y_temp <= 32'b00111100010011111011111000011100;
end
if( x <= 32'b11000000100010110011001100110011 && x > 32'b11000000100010101110000101001000)
begin
	y_temp <= 32'b00111100010100011100110111000001;
end
if( x <= 32'b11000000100010101110000101001000 && x > 32'b11000000100010101000111101011100)
begin
	y_temp <= 32'b00111100010100111110001010010000;
end
if( x <= 32'b11000000100010101000111101011100 && x > 32'b11000000100010100011110101110001)
begin
	y_temp <= 32'b00111100010101011111110010010111;
end
if( x <= 32'b11000000100010100011110101110001 && x > 32'b11000000100010011110101110000101)
begin
	y_temp <= 32'b00111100010110000001101111100010;
end
if( x <= 32'b11000000100010011110101110000101 && x > 32'b11000000100010011001100110011010)
begin
	y_temp <= 32'b00111100010110100100000001111101;
end
if( x <= 32'b11000000100010011001100110011010 && x > 32'b11000000100010010100011110101110)
begin
	y_temp <= 32'b00111100010111000110101001110111;
end
if( x <= 32'b11000000100010010100011110101110 && x > 32'b11000000100010001111010111000011)
begin
	y_temp <= 32'b00111100010111101001100111011011;
end
if( x <= 32'b11000000100010001111010111000011 && x > 32'b11000000100010001010001111010111)
begin
	y_temp <= 32'b00111100011000001100111010110111;
end
if( x <= 32'b11000000100010001010001111010111 && x > 32'b11000000100010000101000111101100)
begin
	y_temp <= 32'b00111100011000110000100100011000;
end
if( x <= 32'b11000000100010000101000111101100 && x > 32'b11000000100010000000000000000000)
begin
	y_temp <= 32'b00111100011001010100100100001011;
end
if( x <= 32'b11000000100010000000000000000000 && x > 32'b11000000100001111010111000010100)
begin
	y_temp <= 32'b00111100011001111000111010011111;
end
if( x <= 32'b11000000100001111010111000010100 && x > 32'b11000000100001110101110000101001)
begin
	y_temp <= 32'b00111100011010011101100111100001;
end
if( x <= 32'b11000000100001110101110000101001 && x > 32'b11000000100001110000101000111101)
begin
	y_temp <= 32'b00111100011011000010101011011110;
end
if( x <= 32'b11000000100001110000101000111101 && x > 32'b11000000100001101011100001010010)
begin
	y_temp <= 32'b00111100011011101000000110100101;
end
if( x <= 32'b11000000100001101011100001010010 && x > 32'b11000000100001100110011001100110)
begin
	y_temp <= 32'b00111100011100001101111001000011;
end
if( x <= 32'b11000000100001100110011001100110 && x > 32'b11000000100001100001010001111011)
begin
	y_temp <= 32'b00111100011100110100000011000111;
end
if( x <= 32'b11000000100001100001010001111011 && x > 32'b11000000100001011100001010001111)
begin
	y_temp <= 32'b00111100011101011010100100111111;
end
if( x <= 32'b11000000100001011100001010001111 && x > 32'b11000000100001010111000010100100)
begin
	y_temp <= 32'b00111100011110000001011110111001;
end
if( x <= 32'b11000000100001010111000010100100 && x > 32'b11000000100001010001111010111000)
begin
	y_temp <= 32'b00111100011110101000110001000100;
end
if( x <= 32'b11000000100001010001111010111000 && x > 32'b11000000100001001100110011001101)
begin
	y_temp <= 32'b00111100011111010000011011101110;
end
if( x <= 32'b11000000100001001100110011001101 && x > 32'b11000000100001000111101011100001)
begin
	y_temp <= 32'b00111100011111111000011111000111;
end
if( x <= 32'b11000000100001000111101011100001 && x > 32'b11000000100001000010100011110110)
begin
	y_temp <= 32'b00111100100000010000011101101110;
end
if( x <= 32'b11000000100001000010100011110110 && x > 32'b11000000100000111101011100001010)
begin
	y_temp <= 32'b00111100100000100100111000011111;
end
if( x <= 32'b11000000100000111101011100001010 && x > 32'b11000000100000111000010100011111)
begin
	y_temp <= 32'b00111100100000111001011111111110;
end
if( x <= 32'b11000000100000111000010100011111 && x > 32'b11000000100000110011001100110011)
begin
	y_temp <= 32'b00111100100001001110010100010001;
end
if( x <= 32'b11000000100000110011001100110011 && x > 32'b11000000100000101110000101001000)
begin
	y_temp <= 32'b00111100100001100011010101100010;
end
if( x <= 32'b11000000100000101110000101001000 && x > 32'b11000000100000101000111101011100)
begin
	y_temp <= 32'b00111100100001111000100011111000;
end
if( x <= 32'b11000000100000101000111101011100 && x > 32'b11000000100000100011110101110001)
begin
	y_temp <= 32'b00111100100010001101111111011010;
end
if( x <= 32'b11000000100000100011110101110001 && x > 32'b11000000100000011110101110000101)
begin
	y_temp <= 32'b00111100100010100011101000010001;
end
if( x <= 32'b11000000100000011110101110000101 && x > 32'b11000000100000011001100110011010)
begin
	y_temp <= 32'b00111100100010111001011110100100;
end
if( x <= 32'b11000000100000011001100110011010 && x > 32'b11000000100000010100011110101110)
begin
	y_temp <= 32'b00111100100011001111100010011100;
end
if( x <= 32'b11000000100000010100011110101110 && x > 32'b11000000100000001111010111000011)
begin
	y_temp <= 32'b00111100100011100101110100000001;
end
if( x <= 32'b11000000100000001111010111000011 && x > 32'b11000000100000001010001111010111)
begin
	y_temp <= 32'b00111100100011111100010011011011;
end
if( x <= 32'b11000000100000001010001111010111 && x > 32'b11000000100000000101000111101100)
begin
	y_temp <= 32'b00111100100100010011000000110010;
end
if( x <= 32'b11000000100000000101000111101100 && x > 32'b11000000100000000000000000000000)
begin
	y_temp <= 32'b00111100100100101001111100001110;
end
if( x <= 32'b11000000100000000000000000000000 && x > 32'b11000000011111110101110000101001)
begin
	y_temp <= 32'b00111100100101000001000101111000;
end
if( x <= 32'b11000000011111110101110000101001 && x > 32'b11000000011111101011100001010010)
begin
	y_temp <= 32'b00111100100101011000011101111001;
end
if( x <= 32'b11000000011111101011100001010010 && x > 32'b11000000011111100001010001111011)
begin
	y_temp <= 32'b00111100100101110000000100011001;
end
if( x <= 32'b11000000011111100001010001111011 && x > 32'b11000000011111010111000010100100)
begin
	y_temp <= 32'b00111100100110000111111001100000;
end
if( x <= 32'b11000000011111010111000010100100 && x > 32'b11000000011111001100110011001101)
begin
	y_temp <= 32'b00111100100110011111111101010111;
end
if( x <= 32'b11000000011111001100110011001101 && x > 32'b11000000011111000010100011110110)
begin
	y_temp <= 32'b00111100100110111000010000001000;
end
if( x <= 32'b11000000011111000010100011110110 && x > 32'b11000000011110111000010100011111)
begin
	y_temp <= 32'b00111100100111010000110001111010;
end
if( x <= 32'b11000000011110111000010100011111 && x > 32'b11000000011110101110000101001000)
begin
	y_temp <= 32'b00111100100111101001100010111000;
end
if( x <= 32'b11000000011110101110000101001000 && x > 32'b11000000011110100011110101110001)
begin
	y_temp <= 32'b00111100101000000010100011001001;
end
if( x <= 32'b11000000011110100011110101110001 && x > 32'b11000000011110011001100110011010)
begin
	y_temp <= 32'b00111100101000011011110010110110;
end
if( x <= 32'b11000000011110011001100110011010 && x > 32'b11000000011110001111010111000011)
begin
	y_temp <= 32'b00111100101000110101010010001010;
end
if( x <= 32'b11000000011110001111010111000011 && x > 32'b11000000011110000101000111101100)
begin
	y_temp <= 32'b00111100101001001111000001001101;
end
if( x <= 32'b11000000011110000101000111101100 && x > 32'b11000000011101111010111000010100)
begin
	y_temp <= 32'b00111100101001101001000000001001;
end
if( x <= 32'b11000000011101111010111000010100 && x > 32'b11000000011101110000101000111101)
begin
	y_temp <= 32'b00111100101010000011001111000111;
end
if( x <= 32'b11000000011101110000101000111101 && x > 32'b11000000011101100110011001100110)
begin
	y_temp <= 32'b00111100101010011101101110010000;
end
if( x <= 32'b11000000011101100110011001100110 && x > 32'b11000000011101011100001010001111)
begin
	y_temp <= 32'b00111100101010111000011101101101;
end
if( x <= 32'b11000000011101011100001010001111 && x > 32'b11000000011101010001111010111000)
begin
	y_temp <= 32'b00111100101011010011011101101010;
end
if( x <= 32'b11000000011101010001111010111000 && x > 32'b11000000011101000111101011100001)
begin
	y_temp <= 32'b00111100101011101110101110001110;
end
if( x <= 32'b11000000011101000111101011100001 && x > 32'b11000000011100111101011100001010)
begin
	y_temp <= 32'b00111100101100001010001111100101;
end
if( x <= 32'b11000000011100111101011100001010 && x > 32'b11000000011100110011001100110011)
begin
	y_temp <= 32'b00111100101100100110000001110111;
end
if( x <= 32'b11000000011100110011001100110011 && x > 32'b11000000011100101000111101011100)
begin
	y_temp <= 32'b00111100101101000010000101001111;
end
if( x <= 32'b11000000011100101000111101011100 && x > 32'b11000000011100011110101110000101)
begin
	y_temp <= 32'b00111100101101011110011001110111;
end
if( x <= 32'b11000000011100011110101110000101 && x > 32'b11000000011100010100011110101110)
begin
	y_temp <= 32'b00111100101101111010111111111001;
end
if( x <= 32'b11000000011100010100011110101110 && x > 32'b11000000011100001010001111010111)
begin
	y_temp <= 32'b00111100101110010111110111011111;
end
if( x <= 32'b11000000011100001010001111010111 && x > 32'b11000000011100000000000000000000)
begin
	y_temp <= 32'b00111100101110110101000000110011;
end
if( x <= 32'b11000000011100000000000000000000 && x > 32'b11000000011011110101110000101001)
begin
	y_temp <= 32'b00111100101111010010011100000000;
end
if( x <= 32'b11000000011011110101110000101001 && x > 32'b11000000011011101011100001010010)
begin
	y_temp <= 32'b00111100101111110000001001010000;
end
if( x <= 32'b11000000011011101011100001010010 && x > 32'b11000000011011100001010001111011)
begin
	y_temp <= 32'b00111100110000001110001000101101;
end
if( x <= 32'b11000000011011100001010001111011 && x > 32'b11000000011011010111000010100100)
begin
	y_temp <= 32'b00111100110000101100011010100011;
end
if( x <= 32'b11000000011011010111000010100100 && x > 32'b11000000011011001100110011001101)
begin
	y_temp <= 32'b00111100110001001010111110111011;
end
if( x <= 32'b11000000011011001100110011001101 && x > 32'b11000000011011000010100011110110)
begin
	y_temp <= 32'b00111100110001101001110110000001;
end
if( x <= 32'b11000000011011000010100011110110 && x > 32'b11000000011010111000010100011111)
begin
	y_temp <= 32'b00111100110010001001000000000000;
end
if( x <= 32'b11000000011010111000010100011111 && x > 32'b11000000011010101110000101001000)
begin
	y_temp <= 32'b00111100110010101000011101000010;
end
if( x <= 32'b11000000011010101110000101001000 && x > 32'b11000000011010100011110101110001)
begin
	y_temp <= 32'b00111100110011001000001101010011;
end
if( x <= 32'b11000000011010100011110101110001 && x > 32'b11000000011010011001100110011010)
begin
	y_temp <= 32'b00111100110011101000010000111101;
end
if( x <= 32'b11000000011010011001100110011010 && x > 32'b11000000011010001111010111000011)
begin
	y_temp <= 32'b00111100110100001000101000001100;
end
if( x <= 32'b11000000011010001111010111000011 && x > 32'b11000000011010000101000111101100)
begin
	y_temp <= 32'b00111100110100101001010011001011;
end
if( x <= 32'b11000000011010000101000111101100 && x > 32'b11000000011001111010111000010100)
begin
	y_temp <= 32'b00111100110101001010010010000110;
end
if( x <= 32'b11000000011001111010111000010100 && x > 32'b11000000011001110000101000111101)
begin
	y_temp <= 32'b00111100110101101011100101001000;
end
if( x <= 32'b11000000011001110000101000111101 && x > 32'b11000000011001100110011001100110)
begin
	y_temp <= 32'b00111100110110001101001100011100;
end
if( x <= 32'b11000000011001100110011001100110 && x > 32'b11000000011001011100001010001111)
begin
	y_temp <= 32'b00111100110110101111001000001110;
end
if( x <= 32'b11000000011001011100001010001111 && x > 32'b11000000011001010001111010111000)
begin
	y_temp <= 32'b00111100110111010001011000101010;
end
if( x <= 32'b11000000011001010001111010111000 && x > 32'b11000000011001000111101011100001)
begin
	y_temp <= 32'b00111100110111110011111101111100;
end
if( x <= 32'b11000000011001000111101011100001 && x > 32'b11000000011000111101011100001010)
begin
	y_temp <= 32'b00111100111000010110111000001111;
end
if( x <= 32'b11000000011000111101011100001010 && x > 32'b11000000011000110011001100110011)
begin
	y_temp <= 32'b00111100111000111010000111110000;
end
if( x <= 32'b11000000011000110011001100110011 && x > 32'b11000000011000101000111101011100)
begin
	y_temp <= 32'b00111100111001011101101100101011;
end
if( x <= 32'b11000000011000101000111101011100 && x > 32'b11000000011000011110101110000101)
begin
	y_temp <= 32'b00111100111010000001100111001100;
end
if( x <= 32'b11000000011000011110101110000101 && x > 32'b11000000011000010100011110101110)
begin
	y_temp <= 32'b00111100111010100101110111011111;
end
if( x <= 32'b11000000011000010100011110101110 && x > 32'b11000000011000001010001111010111)
begin
	y_temp <= 32'b00111100111011001010011101110001;
end
if( x <= 32'b11000000011000001010001111010111 && x > 32'b11000000011000000000000000000000)
begin
	y_temp <= 32'b00111100111011101111011010001110;
end
if( x <= 32'b11000000011000000000000000000000 && x > 32'b11000000010111110101110000101001)
begin
	y_temp <= 32'b00111100111100010100101101000010;
end
if( x <= 32'b11000000010111110101110000101001 && x > 32'b11000000010111101011100001010010)
begin
	y_temp <= 32'b00111100111100111010010110011011;
end
if( x <= 32'b11000000010111101011100001010010 && x > 32'b11000000010111100001010001111011)
begin
	y_temp <= 32'b00111100111101100000010110100101;
end
if( x <= 32'b11000000010111100001010001111011 && x > 32'b11000000010111010111000010100100)
begin
	y_temp <= 32'b00111100111110000110101101101101;
end
if( x <= 32'b11000000010111010111000010100100 && x > 32'b11000000010111001100110011001101)
begin
	y_temp <= 32'b00111100111110101101011100000000;
end
if( x <= 32'b11000000010111001100110011001101 && x > 32'b11000000010111000010100011110110)
begin
	y_temp <= 32'b00111100111111010100100001101011;
end
if( x <= 32'b11000000010111000010100011110110 && x > 32'b11000000010110111000010100011111)
begin
	y_temp <= 32'b00111100111111111011111110111011;
end
if( x <= 32'b11000000010110111000010100011111 && x > 32'b11000000010110101110000101001000)
begin
	y_temp <= 32'b00111101000000010001111001111111;
end
if( x <= 32'b11000000010110101110000101001000 && x > 32'b11000000010110100011110101110001)
begin
	y_temp <= 32'b00111101000000100110000000100000;
end
if( x <= 32'b11000000010110100011110101110001 && x > 32'b11000000010110011001100110011010)
begin
	y_temp <= 32'b00111101000000111010010011000111;
end
if( x <= 32'b11000000010110011001100110011010 && x > 32'b11000000010110001111010111000011)
begin
	y_temp <= 32'b00111101000001001110110001111100;
end
if( x <= 32'b11000000010110001111010111000011 && x > 32'b11000000010110000101000111101100)
begin
	y_temp <= 32'b00111101000001100011011101000110;
end
if( x <= 32'b11000000010110000101000111101100 && x > 32'b11000000010101111010111000010100)
begin
	y_temp <= 32'b00111101000001111000010100101010;
end
if( x <= 32'b11000000010101111010111000010100 && x > 32'b11000000010101110000101000111101)
begin
	y_temp <= 32'b00111101000010001101011000110000;
end
if( x <= 32'b11000000010101110000101000111101 && x > 32'b11000000010101100110011001100110)
begin
	y_temp <= 32'b00111101000010100010101001011111;
end
if( x <= 32'b11000000010101100110011001100110 && x > 32'b11000000010101011100001010001111)
begin
	y_temp <= 32'b00111101000010111000000110111110;
end
if( x <= 32'b11000000010101011100001010001111 && x > 32'b11000000010101010001111010111000)
begin
	y_temp <= 32'b00111101000011001101110001010100;
end
if( x <= 32'b11000000010101010001111010111000 && x > 32'b11000000010101000111101011100001)
begin
	y_temp <= 32'b00111101000011100011101000101000;
end
if( x <= 32'b11000000010101000111101011100001 && x > 32'b11000000010100111101011100001010)
begin
	y_temp <= 32'b00111101000011111001101101000001;
end
if( x <= 32'b11000000010100111101011100001010 && x > 32'b11000000010100110011001100110011)
begin
	y_temp <= 32'b00111101000100001111111110100111;
end
if( x <= 32'b11000000010100110011001100110011 && x > 32'b11000000010100101000111101011100)
begin
	y_temp <= 32'b00111101000100100110011101100000;
end
if( x <= 32'b11000000010100101000111101011100 && x > 32'b11000000010100011110101110000101)
begin
	y_temp <= 32'b00111101000100111101001001110101;
end
if( x <= 32'b11000000010100011110101110000101 && x > 32'b11000000010100010100011110101110)
begin
	y_temp <= 32'b00111101000101010100000011101011;
end
if( x <= 32'b11000000010100010100011110101110 && x > 32'b11000000010100001010001111010111)
begin
	y_temp <= 32'b00111101000101101011001011001100;
end
if( x <= 32'b11000000010100001010001111010111 && x > 32'b11000000010100000000000000000000)
begin
	y_temp <= 32'b00111101000110000010100000011110;
end
if( x <= 32'b11000000010100000000000000000000 && x > 32'b11000000010011110101110000101001)
begin
	y_temp <= 32'b00111101000110011010000011101001;
end
if( x <= 32'b11000000010011110101110000101001 && x > 32'b11000000010011101011100001010010)
begin
	y_temp <= 32'b00111101000110110001110100110100;
end
if( x <= 32'b11000000010011101011100001010010 && x > 32'b11000000010011100001010001111011)
begin
	y_temp <= 32'b00111101000111001001110100000111;
end
if( x <= 32'b11000000010011100001010001111011 && x > 32'b11000000010011010111000010100100)
begin
	y_temp <= 32'b00111101000111100010000001101010;
end
if( x <= 32'b11000000010011010111000010100100 && x > 32'b11000000010011001100110011001101)
begin
	y_temp <= 32'b00111101000111111010011101100100;
end
if( x <= 32'b11000000010011001100110011001101 && x > 32'b11000000010011000010100011110110)
begin
	y_temp <= 32'b00111101001000010011000111111110;
end
if( x <= 32'b11000000010011000010100011110110 && x > 32'b11000000010010111000010100011111)
begin
	y_temp <= 32'b00111101001000101100000000111110;
end
if( x <= 32'b11000000010010111000010100011111 && x > 32'b11000000010010101110000101001000)
begin
	y_temp <= 32'b00111101001001000101001000101101;
end
if( x <= 32'b11000000010010101110000101001000 && x > 32'b11000000010010100011110101110001)
begin
	y_temp <= 32'b00111101001001011110011111010011;
end
if( x <= 32'b11000000010010100011110101110001 && x > 32'b11000000010010011001100110011010)
begin
	y_temp <= 32'b00111101001001111000000100111000;
end
if( x <= 32'b11000000010010011001100110011010 && x > 32'b11000000010010001111010111000011)
begin
	y_temp <= 32'b00111101001010010001111001100011;
end
if( x <= 32'b11000000010010001111010111000011 && x > 32'b11000000010010000101000111101100)
begin
	y_temp <= 32'b00111101001010101011111101011101;
end
if( x <= 32'b11000000010010000101000111101100 && x > 32'b11000000010001111010111000010100)
begin
	y_temp <= 32'b00111101001011000110010000101110;
end
if( x <= 32'b11000000010001111010111000010100 && x > 32'b11000000010001110000101000111101)
begin
	y_temp <= 32'b00111101001011100000110011011111;
end
if( x <= 32'b11000000010001110000101000111101 && x > 32'b11000000010001100110011001100110)
begin
	y_temp <= 32'b00111101001011111011100101110110;
end
if( x <= 32'b11000000010001100110011001100110 && x > 32'b11000000010001011100001010001111)
begin
	y_temp <= 32'b00111101001100010110100111111110;
end
if( x <= 32'b11000000010001011100001010001111 && x > 32'b11000000010001010001111010111000)
begin
	y_temp <= 32'b00111101001100110001111001111101;
end
if( x <= 32'b11000000010001010001111010111000 && x > 32'b11000000010001000111101011100001)
begin
	y_temp <= 32'b00111101001101001101011011111101;
end
if( x <= 32'b11000000010001000111101011100001 && x > 32'b11000000010000111101011100001010)
begin
	y_temp <= 32'b00111101001101101001001110000101;
end
if( x <= 32'b11000000010000111101011100001010 && x > 32'b11000000010000110011001100110011)
begin
	y_temp <= 32'b00111101001110000101010000011111;
end
if( x <= 32'b11000000010000110011001100110011 && x > 32'b11000000010000101000111101011100)
begin
	y_temp <= 32'b00111101001110100001100011010011;
end
if( x <= 32'b11000000010000101000111101011100 && x > 32'b11000000010000011110101110000101)
begin
	y_temp <= 32'b00111101001110111110000110101001;
end
if( x <= 32'b11000000010000011110101110000101 && x > 32'b11000000010000010100011110101110)
begin
	y_temp <= 32'b00111101001111011010111010101010;
end
if( x <= 32'b11000000010000010100011110101110 && x > 32'b11000000010000001010001111010111)
begin
	y_temp <= 32'b00111101001111110111111111011111;
end
if( x <= 32'b11000000010000001010001111010111 && x > 32'b11000000010000000000000000000000)
begin
	y_temp <= 32'b00111101010000010101010101010000;
end
if( x <= 32'b11000000010000000000000000000000 && x > 32'b11000000001111110101110000101001)
begin
	y_temp <= 32'b00111101010000110010111100000110;
end
if( x <= 32'b11000000001111110101110000101001 && x > 32'b11000000001111101011100001010010)
begin
	y_temp <= 32'b00111101010001010000110100001011;
end
if( x <= 32'b11000000001111101011100001010010 && x > 32'b11000000001111100001010001111011)
begin
	y_temp <= 32'b00111101010001101110111101100111;
end
if( x <= 32'b11000000001111100001010001111011 && x > 32'b11000000001111010111000010100100)
begin
	y_temp <= 32'b00111101010010001101011000100010;
end
if( x <= 32'b11000000001111010111000010100100 && x > 32'b11000000001111001100110011001101)
begin
	y_temp <= 32'b00111101010010101100000101000111;
end
if( x <= 32'b11000000001111001100110011001101 && x > 32'b11000000001111000010100011110110)
begin
	y_temp <= 32'b00111101010011001011000011011101;
end
if( x <= 32'b11000000001111000010100011110110 && x > 32'b11000000001110111000010100011111)
begin
	y_temp <= 32'b00111101010011101010010011101111;
end
if( x <= 32'b11000000001110111000010100011111 && x > 32'b11000000001110101110000101001000)
begin
	y_temp <= 32'b00111101010100001001110110000100;
end
if( x <= 32'b11000000001110101110000101001000 && x > 32'b11000000001110100011110101110001)
begin
	y_temp <= 32'b00111101010100101001101010101000;
end
if( x <= 32'b11000000001110100011110101110001 && x > 32'b11000000001110011001100110011010)
begin
	y_temp <= 32'b00111101010101001001110001100001;
end
if( x <= 32'b11000000001110011001100110011010 && x > 32'b11000000001110001111010111000011)
begin
	y_temp <= 32'b00111101010101101010001010111011;
end
if( x <= 32'b11000000001110001111010111000011 && x > 32'b11000000001110000101000111101100)
begin
	y_temp <= 32'b00111101010110001010110110111110;
end
if( x <= 32'b11000000001110000101000111101100 && x > 32'b11000000001101111010111000010100)
begin
	y_temp <= 32'b00111101010110101011110101110011;
end
if( x <= 32'b11000000001101111010111000010100 && x > 32'b11000000001101110000101000111101)
begin
	y_temp <= 32'b00111101010111001101000111100101;
end
if( x <= 32'b11000000001101110000101000111101 && x > 32'b11000000001101100110011001100110)
begin
	y_temp <= 32'b00111101010111101110101100011100;
end
if( x <= 32'b11000000001101100110011001100110 && x > 32'b11000000001101011100001010001111)
begin
	y_temp <= 32'b00111101011000010000100100100010;
end
if( x <= 32'b11000000001101011100001010001111 && x > 32'b11000000001101010001111010111000)
begin
	y_temp <= 32'b00111101011000110010110000000001;
end
if( x <= 32'b11000000001101010001111010111000 && x > 32'b11000000001101000111101011100001)
begin
	y_temp <= 32'b00111101011001010101001111000010;
end
if( x <= 32'b11000000001101000111101011100001 && x > 32'b11000000001100111101011100001010)
begin
	y_temp <= 32'b00111101011001111000000001101110;
end
if( x <= 32'b11000000001100111101011100001010 && x > 32'b11000000001100110011001100110011)
begin
	y_temp <= 32'b00111101011010011011001000010001;
end
if( x <= 32'b11000000001100110011001100110011 && x > 32'b11000000001100101000111101011100)
begin
	y_temp <= 32'b00111101011010111110100010110011;
end
if( x <= 32'b11000000001100101000111101011100 && x > 32'b11000000001100011110101110000101)
begin
	y_temp <= 32'b00111101011011100010010001011110;
end
if( x <= 32'b11000000001100011110101110000101 && x > 32'b11000000001100010100011110101110)
begin
	y_temp <= 32'b00111101011100000110010100011100;
end
if( x <= 32'b11000000001100010100011110101110 && x > 32'b11000000001100001010001111010111)
begin
	y_temp <= 32'b00111101011100101010101011110111;
end
if( x <= 32'b11000000001100001010001111010111 && x > 32'b11000000001100000000000000000000)
begin
	y_temp <= 32'b00111101011101001111010111111001;
end
if( x <= 32'b11000000001100000000000000000000 && x > 32'b11000000001011110101110000101001)
begin
	y_temp <= 32'b00111101011101110100011000101011;
end
if( x <= 32'b11000000001011110101110000101001 && x > 32'b11000000001011101011100001010010)
begin
	y_temp <= 32'b00111101011110011001101110011001;
end
if( x <= 32'b11000000001011101011100001010010 && x > 32'b11000000001011100001010001111011)
begin
	y_temp <= 32'b00111101011110111111011001001011;
end
if( x <= 32'b11000000001011100001010001111011 && x > 32'b11000000001011010111000010100100)
begin
	y_temp <= 32'b00111101011111100101011001001101;
end
if( x <= 32'b11000000001011010111000010100100 && x > 32'b11000000001011001100110011001101)
begin
	y_temp <= 32'b00111101100000000101110111010100;
end
if( x <= 32'b11000000001011001100110011001101 && x > 32'b11000000001011000010100011110110)
begin
	y_temp <= 32'b00111101100000011001001100110011;
end
if( x <= 32'b11000000001011000010100011110110 && x > 32'b11000000001010111000010100011111)
begin
	y_temp <= 32'b00111101100000101100101101001001;
end
if( x <= 32'b11000000001010111000010100011111 && x > 32'b11000000001010101110000101001000)
begin
	y_temp <= 32'b00111101100001000000011000011010;
end
if( x <= 32'b11000000001010101110000101001000 && x > 32'b11000000001010100011110101110001)
begin
	y_temp <= 32'b00111101100001010100001110101101;
end
if( x <= 32'b11000000001010100011110101110001 && x > 32'b11000000001010011001100110011010)
begin
	y_temp <= 32'b00111101100001101000010000000110;
end
if( x <= 32'b11000000001010011001100110011010 && x > 32'b11000000001010001111010111000011)
begin
	y_temp <= 32'b00111101100001111100011100101011;
end
if( x <= 32'b11000000001010001111010111000011 && x > 32'b11000000001010000101000111101100)
begin
	y_temp <= 32'b00111101100010010000110100100000;
end
if( x <= 32'b11000000001010000101000111101100 && x > 32'b11000000001001111010111000010100)
begin
	y_temp <= 32'b00111101100010100101010111101011;
end
if( x <= 32'b11000000001001111010111000010100 && x > 32'b11000000001001110000101000111101)
begin
	y_temp <= 32'b00111101100010111010000110010010;
end
if( x <= 32'b11000000001001110000101000111101 && x > 32'b11000000001001100110011001100110)
begin
	y_temp <= 32'b00111101100011001111000000011001;
end
if( x <= 32'b11000000001001100110011001100110 && x > 32'b11000000001001011100001010001111)
begin
	y_temp <= 32'b00111101100011100100000110000101;
end
if( x <= 32'b11000000001001011100001010001111 && x > 32'b11000000001001010001111010111000)
begin
	y_temp <= 32'b00111101100011111001010111011100;
end
if( x <= 32'b11000000001001010001111010111000 && x > 32'b11000000001001000111101011100001)
begin
	y_temp <= 32'b00111101100100001110110100100100;
end
if( x <= 32'b11000000001001000111101011100001 && x > 32'b11000000001000111101011100001010)
begin
	y_temp <= 32'b00111101100100100100011101100010;
end
if( x <= 32'b11000000001000111101011100001010 && x > 32'b11000000001000110011001100110011)
begin
	y_temp <= 32'b00111101100100111010010010011010;
end
if( x <= 32'b11000000001000110011001100110011 && x > 32'b11000000001000101000111101011100)
begin
	y_temp <= 32'b00111101100101010000010011010011;
end
if( x <= 32'b11000000001000101000111101011100 && x > 32'b11000000001000011110101110000101)
begin
	y_temp <= 32'b00111101100101100110100000010010;
end
if( x <= 32'b11000000001000011110101110000101 && x > 32'b11000000001000010100011110101110)
begin
	y_temp <= 32'b00111101100101111100111001011100;
end
if( x <= 32'b11000000001000010100011110101110 && x > 32'b11000000001000001010001111010111)
begin
	y_temp <= 32'b00111101100110010011011110110110;
end
if( x <= 32'b11000000001000001010001111010111 && x > 32'b11000000001000000000000000000000)
begin
	y_temp <= 32'b00111101100110101010010000100110;
end
if( x <= 32'b11000000001000000000000000000000 && x > 32'b11000000000111110101110000101001)
begin
	y_temp <= 32'b00111101100111000001001110110010;
end
if( x <= 32'b11000000000111110101110000101001 && x > 32'b11000000000111101011100001010010)
begin
	y_temp <= 32'b00111101100111011000011001011111;
end
if( x <= 32'b11000000000111101011100001010010 && x > 32'b11000000000111100001010001111011)
begin
	y_temp <= 32'b00111101100111101111110000110010;
end
if( x <= 32'b11000000000111100001010001111011 && x > 32'b11000000000111010111000010100100)
begin
	y_temp <= 32'b00111101101000000111010100110001;
end
if( x <= 32'b11000000000111010111000010100100 && x > 32'b11000000000111001100110011001101)
begin
	y_temp <= 32'b00111101101000011111000101100001;
end
if( x <= 32'b11000000000111001100110011001101 && x > 32'b11000000000111000010100011110110)
begin
	y_temp <= 32'b00111101101000110111000011001000;
end
if( x <= 32'b11000000000111000010100011110110 && x > 32'b11000000000110111000010100011111)
begin
	y_temp <= 32'b00111101101001001111001101101100;
end
if( x <= 32'b11000000000110111000010100011111 && x > 32'b11000000000110101110000101001000)
begin
	y_temp <= 32'b00111101101001100111100101010001;
end
if( x <= 32'b11000000000110101110000101001000 && x > 32'b11000000000110100011110101110001)
begin
	y_temp <= 32'b00111101101010000000001001111110;
end
if( x <= 32'b11000000000110100011110101110001 && x > 32'b11000000000110011001100110011010)
begin
	y_temp <= 32'b00111101101010011000111011110111;
end
if( x <= 32'b11000000000110011001100110011010 && x > 32'b11000000000110001111010111000011)
begin
	y_temp <= 32'b00111101101010110001111011000011;
end
if( x <= 32'b11000000000110001111010111000011 && x > 32'b11000000000110000101000111101100)
begin
	y_temp <= 32'b00111101101011001011000111100111;
end
if( x <= 32'b11000000000110000101000111101100 && x > 32'b11000000000101111010111000010100)
begin
	y_temp <= 32'b00111101101011100100100001101000;
end
if( x <= 32'b11000000000101111010111000010100 && x > 32'b11000000000101110000101000111101)
begin
	y_temp <= 32'b00111101101011111110001001001101;
end
if( x <= 32'b11000000000101110000101000111101 && x > 32'b11000000000101100110011001100110)
begin
	y_temp <= 32'b00111101101100010111111110011010;
end
if( x <= 32'b11000000000101100110011001100110 && x > 32'b11000000000101011100001010001111)
begin
	y_temp <= 32'b00111101101100110010000001010110;
end
if( x <= 32'b11000000000101011100001010001111 && x > 32'b11000000000101010001111010111000)
begin
	y_temp <= 32'b00111101101101001100010010000110;
end
if( x <= 32'b11000000000101010001111010111000 && x > 32'b11000000000101000111101011100001)
begin
	y_temp <= 32'b00111101101101100110110000101111;
end
if( x <= 32'b11000000000101000111101011100001 && x > 32'b11000000000100111101011100001010)
begin
	y_temp <= 32'b00111101101110000001011101010110;
end
if( x <= 32'b11000000000100111101011100001010 && x > 32'b11000000000100110011001100110011)
begin
	y_temp <= 32'b00111101101110011100011000000011;
end
if( x <= 32'b11000000000100110011001100110011 && x > 32'b11000000000100101000111101011100)
begin
	y_temp <= 32'b00111101101110110111100000111010;
end
if( x <= 32'b11000000000100101000111101011100 && x > 32'b11000000000100011110101110000101)
begin
	y_temp <= 32'b00111101101111010010111000000000;
end
if( x <= 32'b11000000000100011110101110000101 && x > 32'b11000000000100010100011110101110)
begin
	y_temp <= 32'b00111101101111101110011101011100;
end
if( x <= 32'b11000000000100010100011110101110 && x > 32'b11000000000100001010001111010111)
begin
	y_temp <= 32'b00111101110000001010010001010011;
end
if( x <= 32'b11000000000100001010001111010111 && x > 32'b11000000000100000000000000000000)
begin
	y_temp <= 32'b00111101110000100110010011101011;
end
if( x <= 32'b11000000000100000000000000000000 && x > 32'b11000000000011110101110000101001)
begin
	y_temp <= 32'b00111101110001000010100100101001;
end
if( x <= 32'b11000000000011110101110000101001 && x > 32'b11000000000011101011100001010010)
begin
	y_temp <= 32'b00111101110001011111000100010010;
end
if( x <= 32'b11000000000011101011100001010010 && x > 32'b11000000000011100001010001111011)
begin
	y_temp <= 32'b00111101110001111011110010101101;
end
if( x <= 32'b11000000000011100001010001111011 && x > 32'b11000000000011010111000010100100)
begin
	y_temp <= 32'b00111101110010011000101111111110;
end
if( x <= 32'b11000000000011010111000010100100 && x > 32'b11000000000011001100110011001101)
begin
	y_temp <= 32'b00111101110010110101111100001101;
end
if( x <= 32'b11000000000011001100110011001101 && x > 32'b11000000000011000010100011110110)
begin
	y_temp <= 32'b00111101110011010011010111011101;
end
if( x <= 32'b11000000000011000010100011110110 && x > 32'b11000000000010111000010100011111)
begin
	y_temp <= 32'b00111101110011110001000001110101;
end
if( x <= 32'b11000000000010111000010100011111 && x > 32'b11000000000010101110000101001000)
begin
	y_temp <= 32'b00111101110100001110111011011001;
end
if( x <= 32'b11000000000010101110000101001000 && x > 32'b11000000000010100011110101110001)
begin
	y_temp <= 32'b00111101110100101101000100010001;
end
if( x <= 32'b11000000000010100011110101110001 && x > 32'b11000000000010011001100110011010)
begin
	y_temp <= 32'b00111101110101001011011100100001;
end
if( x <= 32'b11000000000010011001100110011010 && x > 32'b11000000000010001111010111000011)
begin
	y_temp <= 32'b00111101110101101010000100001111;
end
if( x <= 32'b11000000000010001111010111000011 && x > 32'b11000000000010000101000111101100)
begin
	y_temp <= 32'b00111101110110001000111011011111;
end
if( x <= 32'b11000000000010000101000111101100 && x > 32'b11000000000001111010111000010100)
begin
	y_temp <= 32'b00111101110110101000000010011001;
end
if( x <= 32'b11000000000001111010111000010100 && x > 32'b11000000000001110000101000111101)
begin
	y_temp <= 32'b00111101110111000111011001000001;
end
if( x <= 32'b11000000000001110000101000111101 && x > 32'b11000000000001100110011001100110)
begin
	y_temp <= 32'b00111101110111100110111111011101;
end
if( x <= 32'b11000000000001100110011001100110 && x > 32'b11000000000001011100001010001111)
begin
	y_temp <= 32'b00111101111000000110110101110001;
end
if( x <= 32'b11000000000001011100001010001111 && x > 32'b11000000000001010001111010111000)
begin
	y_temp <= 32'b00111101111000100110111100000101;
end
if( x <= 32'b11000000000001010001111010111000 && x > 32'b11000000000001000111101011100001)
begin
	y_temp <= 32'b00111101111001000111010010011100;
end
if( x <= 32'b11000000000001000111101011100001 && x > 32'b11000000000000111101011100001010)
begin
	y_temp <= 32'b00111101111001100111111000111101;
end
if( x <= 32'b11000000000000111101011100001010 && x > 32'b11000000000000110011001100110011)
begin
	y_temp <= 32'b00111101111010001000101111101100;
end
if( x <= 32'b11000000000000110011001100110011 && x > 32'b11000000000000101000111101011100)
begin
	y_temp <= 32'b00111101111010101001110110110000;
end
if( x <= 32'b11000000000000101000111101011100 && x > 32'b11000000000000011110101110000101)
begin
	y_temp <= 32'b00111101111011001011001110001110;
end
if( x <= 32'b11000000000000011110101110000101 && x > 32'b11000000000000010100011110101110)
begin
	y_temp <= 32'b00111101111011101100110110001010;
end
if( x <= 32'b11000000000000010100011110101110 && x > 32'b11000000000000001010001111010111)
begin
	y_temp <= 32'b00111101111100001110101110101010;
end
if( x <= 32'b11000000000000001010001111010111 && x > 32'b11000000000000000000000000000000)
begin
	y_temp <= 32'b00111101111100110000110111110011;
end
if( x <= 32'b11000000000000000000000000000000 && x > 32'b10111111111111101011100001010010)
begin
	y_temp <= 32'b00111101111101010011010001101100;
end
if( x <= 32'b10111111111111101011100001010010 && x > 32'b10111111111111010111000010100100)
begin
	y_temp <= 32'b00111101111101110101111100011000;
end
if( x <= 32'b10111111111111010111000010100100 && x > 32'b10111111111111000010100011110110)
begin
	y_temp <= 32'b00111101111110011000110111111101;
end
if( x <= 32'b10111111111111000010100011110110 && x > 32'b10111111111110101110000101001000)
begin
	y_temp <= 32'b00111101111110111100000100100000;
end
if( x <= 32'b10111111111110101110000101001000 && x > 32'b10111111111110011001100110011010)
begin
	y_temp <= 32'b00111101111111011111100010000111;
end
if( x <= 32'b10111111111110011001100110011010 && x > 32'b10111111111110000101000111101100)
begin
	y_temp <= 32'b00111110000000000001101000011011;
end
if( x <= 32'b10111111111110000101000111101100 && x > 32'b10111111111101110000101000111101)
begin
	y_temp <= 32'b00111110000000010011101000011001;
end
if( x <= 32'b10111111111101110000101000111101 && x > 32'b10111111111101011100001010001111)
begin
	y_temp <= 32'b00111110000000100101110001000000;
end
if( x <= 32'b10111111111101011100001010001111 && x > 32'b10111111111101000111101011100001)
begin
	y_temp <= 32'b00111110000000111000000010010100;
end
if( x <= 32'b10111111111101000111101011100001 && x > 32'b10111111111100110011001100110011)
begin
	y_temp <= 32'b00111110000001001010011100010101;
end
if( x <= 32'b10111111111100110011001100110011 && x > 32'b10111111111100011110101110000101)
begin
	y_temp <= 32'b00111110000001011100111111000111;
end
if( x <= 32'b10111111111100011110101110000101 && x > 32'b10111111111100001010001111010111)
begin
	y_temp <= 32'b00111110000001101111101010101100;
end
if( x <= 32'b10111111111100001010001111010111 && x > 32'b10111111111011110101110000101001)
begin
	y_temp <= 32'b00111110000010000010011111000111;
end
if( x <= 32'b10111111111011110101110000101001 && x > 32'b10111111111011100001010001111011)
begin
	y_temp <= 32'b00111110000010010101011100011010;
end
if( x <= 32'b10111111111011100001010001111011 && x > 32'b10111111111011001100110011001101)
begin
	y_temp <= 32'b00111110000010101000100010100111;
end
if( x <= 32'b10111111111011001100110011001101 && x > 32'b10111111111010111000010100011111)
begin
	y_temp <= 32'b00111110000010111011110001110000;
end
if( x <= 32'b10111111111010111000010100011111 && x > 32'b10111111111010100011110101110001)
begin
	y_temp <= 32'b00111110000011001111001001111001;
end
if( x <= 32'b10111111111010100011110101110001 && x > 32'b10111111111010001111010111000011)
begin
	y_temp <= 32'b00111110000011100010101011000011;
end
if( x <= 32'b10111111111010001111010111000011 && x > 32'b10111111111001111010111000010100)
begin
	y_temp <= 32'b00111110000011110110010101010000;
end
if( x <= 32'b10111111111001111010111000010100 && x > 32'b10111111111001100110011001100110)
begin
	y_temp <= 32'b00111110000100001010001000100011;
end
if( x <= 32'b10111111111001100110011001100110 && x > 32'b10111111111001010001111010111000)
begin
	y_temp <= 32'b00111110000100011110000100111111;
end
if( x <= 32'b10111111111001010001111010111000 && x > 32'b10111111111000111101011100001010)
begin
	y_temp <= 32'b00111110000100110010001010100100;
end
if( x <= 32'b10111111111000111101011100001010 && x > 32'b10111111111000101000111101011100)
begin
	y_temp <= 32'b00111110000101000110011001010110;
end
if( x <= 32'b10111111111000101000111101011100 && x > 32'b10111111111000010100011110101110)
begin
	y_temp <= 32'b00111110000101011010110001010111;
end
if( x <= 32'b10111111111000010100011110101110 && x > 32'b10111111111000000000000000000000)
begin
	y_temp <= 32'b00111110000101101111010010101000;
end
if( x <= 32'b10111111111000000000000000000000 && x > 32'b10111111110111101011100001010010)
begin
	y_temp <= 32'b00111110000110000011111101001100;
end
if( x <= 32'b10111111110111101011100001010010 && x > 32'b10111111110111010111000010100100)
begin
	y_temp <= 32'b00111110000110011000110001000101;
end
if( x <= 32'b10111111110111010111000010100100 && x > 32'b10111111110111000010100011110110)
begin
	y_temp <= 32'b00111110000110101101101110010100;
end
if( x <= 32'b10111111110111000010100011110110 && x > 32'b10111111110110101110000101001000)
begin
	y_temp <= 32'b00111110000111000010110100111101;
end
if( x <= 32'b10111111110110101110000101001000 && x > 32'b10111111110110011001100110011010)
begin
	y_temp <= 32'b00111110000111011000000101000000;
end
if( x <= 32'b10111111110110011001100110011010 && x > 32'b10111111110110000101000111101100)
begin
	y_temp <= 32'b00111110000111101101011110100000;
end
if( x <= 32'b10111111110110000101000111101100 && x > 32'b10111111110101110000101000111101)
begin
	y_temp <= 32'b00111110001000000011000001011111;
end
if( x <= 32'b10111111110101110000101000111101 && x > 32'b10111111110101011100001010001111)
begin
	y_temp <= 32'b00111110001000011000101101111110;
end
if( x <= 32'b10111111110101011100001010001111 && x > 32'b10111111110101000111101011100001)
begin
	y_temp <= 32'b00111110001000101110100100000000;
end
if( x <= 32'b10111111110101000111101011100001 && x > 32'b10111111110100110011001100110011)
begin
	y_temp <= 32'b00111110001001000100100011100110;
end
if( x <= 32'b10111111110100110011001100110011 && x > 32'b10111111110100011110101110000101)
begin
	y_temp <= 32'b00111110001001011010101100110001;
end
if( x <= 32'b10111111110100011110101110000101 && x > 32'b10111111110100001010001111010111)
begin
	y_temp <= 32'b00111110001001110000111111100100;
end
if( x <= 32'b10111111110100001010001111010111 && x > 32'b10111111110011110101110000101001)
begin
	y_temp <= 32'b00111110001010000111011100000001;
end
if( x <= 32'b10111111110011110101110000101001 && x > 32'b10111111110011100001010001111011)
begin
	y_temp <= 32'b00111110001010011110000010001000;
end
if( x <= 32'b10111111110011100001010001111011 && x > 32'b10111111110011001100110011001101)
begin
	y_temp <= 32'b00111110001010110100110001111100;
end
if( x <= 32'b10111111110011001100110011001101 && x > 32'b10111111110010111000010100011111)
begin
	y_temp <= 32'b00111110001011001011101011011110;
end
if( x <= 32'b10111111110010111000010100011111 && x > 32'b10111111110010100011110101110001)
begin
	y_temp <= 32'b00111110001011100010101110110000;
end
if( x <= 32'b10111111110010100011110101110001 && x > 32'b10111111110010001111010111000011)
begin
	y_temp <= 32'b00111110001011111001111011110010;
end
if( x <= 32'b10111111110010001111010111000011 && x > 32'b10111111110001111010111000010100)
begin
	y_temp <= 32'b00111110001100010001010010100111;
end
if( x <= 32'b10111111110001111010111000010100 && x > 32'b10111111110001100110011001100110)
begin
	y_temp <= 32'b00111110001100101000110011010000;
end
if( x <= 32'b10111111110001100110011001100110 && x > 32'b10111111110001010001111010111000)
begin
	y_temp <= 32'b00111110001101000000011101101110;
end
if( x <= 32'b10111111110001010001111010111000 && x > 32'b10111111110000111101011100001010)
begin
	y_temp <= 32'b00111110001101011000010010000011;
end
if( x <= 32'b10111111110000111101011100001010 && x > 32'b10111111110000101000111101011100)
begin
	y_temp <= 32'b00111110001101110000010000001111;
end
if( x <= 32'b10111111110000101000111101011100 && x > 32'b10111111110000010100011110101110)
begin
	y_temp <= 32'b00111110001110001000011000010101;
end
if( x <= 32'b10111111110000010100011110101110 && x > 32'b10111111110000000000000000000000)
begin
	y_temp <= 32'b00111110001110100000101010010100;
end
if( x <= 32'b10111111110000000000000000000000 && x > 32'b10111111101111101011100001010010)
begin
	y_temp <= 32'b00111110001110111001000110001110;
end
if( x <= 32'b10111111101111101011100001010010 && x > 32'b10111111101111010111000010100100)
begin
	y_temp <= 32'b00111110001111010001101100000101;
end
if( x <= 32'b10111111101111010111000010100100 && x > 32'b10111111101111000010100011110110)
begin
	y_temp <= 32'b00111110001111101010011011111001;
end
if( x <= 32'b10111111101111000010100011110110 && x > 32'b10111111101110101110000101001000)
begin
	y_temp <= 32'b00111110010000000011010101101011;
end
if( x <= 32'b10111111101110101110000101001000 && x > 32'b10111111101110011001100110011010)
begin
	y_temp <= 32'b00111110010000011100011001011101;
end
if( x <= 32'b10111111101110011001100110011010 && x > 32'b10111111101110000101000111101100)
begin
	y_temp <= 32'b00111110010000110101100111001110;
end
if( x <= 32'b10111111101110000101000111101100 && x > 32'b10111111101101110000101000111101)
begin
	y_temp <= 32'b00111110010001001110111111000000;
end
if( x <= 32'b10111111101101110000101000111101 && x > 32'b10111111101101011100001010001111)
begin
	y_temp <= 32'b00111110010001101000100000110011;
end
if( x <= 32'b10111111101101011100001010001111 && x > 32'b10111111101101000111101011100001)
begin
	y_temp <= 32'b00111110010010000010001100101001;
end
if( x <= 32'b10111111101101000111101011100001 && x > 32'b10111111101100110011001100110011)
begin
	y_temp <= 32'b00111110010010011100000010100001;
end
if( x <= 32'b10111111101100110011001100110011 && x > 32'b10111111101100011110101110000101)
begin
	y_temp <= 32'b00111110010010110110000010011101;
end
if( x <= 32'b10111111101100011110101110000101 && x > 32'b10111111101100001010001111010111)
begin
	y_temp <= 32'b00111110010011010000001100011100;
end
if( x <= 32'b10111111101100001010001111010111 && x > 32'b10111111101011110101110000101001)
begin
	y_temp <= 32'b00111110010011101010100000100000;
end
if( x <= 32'b10111111101011110101110000101001 && x > 32'b10111111101011100001010001111011)
begin
	y_temp <= 32'b00111110010100000100111110101001;
end
if( x <= 32'b10111111101011100001010001111011 && x > 32'b10111111101011001100110011001101)
begin
	y_temp <= 32'b00111110010100011111100110110110;
end
if( x <= 32'b10111111101011001100110011001101 && x > 32'b10111111101010111000010100011111)
begin
	y_temp <= 32'b00111110010100111010011001001001;
end
if( x <= 32'b10111111101010111000010100011111 && x > 32'b10111111101010100011110101110001)
begin
	y_temp <= 32'b00111110010101010101010101100001;
end
if( x <= 32'b10111111101010100011110101110001 && x > 32'b10111111101010001111010111000011)
begin
	y_temp <= 32'b00111110010101110000011011111111;
end
if( x <= 32'b10111111101010001111010111000011 && x > 32'b10111111101001111010111000010100)
begin
	y_temp <= 32'b00111110010110001011101100100011;
end
if( x <= 32'b10111111101001111010111000010100 && x > 32'b10111111101001100110011001100110)
begin
	y_temp <= 32'b00111110010110100111000111001100;
end
if( x <= 32'b10111111101001100110011001100110 && x > 32'b10111111101001010001111010111000)
begin
	y_temp <= 32'b00111110010111000010101011111011;
end
if( x <= 32'b10111111101001010001111010111000 && x > 32'b10111111101000111101011100001010)
begin
	y_temp <= 32'b00111110010111011110011010110000;
end
if( x <= 32'b10111111101000111101011100001010 && x > 32'b10111111101000101000111101011100)
begin
	y_temp <= 32'b00111110010111111010010011101010;
end
if( x <= 32'b10111111101000101000111101011100 && x > 32'b10111111101000010100011110101110)
begin
	y_temp <= 32'b00111110011000010110010110101001;
end
if( x <= 32'b10111111101000010100011110101110 && x > 32'b10111111101000000000000000000000)
begin
	y_temp <= 32'b00111110011000110010100011101110;
end
if( x <= 32'b10111111101000000000000000000000 && x > 32'b10111111100111101011100001010010)
begin
	y_temp <= 32'b00111110011001001110111010110110;
end
if( x <= 32'b10111111100111101011100001010010 && x > 32'b10111111100111010111000010100100)
begin
	y_temp <= 32'b00111110011001101011011100000011;
end
if( x <= 32'b10111111100111010111000010100100 && x > 32'b10111111100111000010100011110110)
begin
	y_temp <= 32'b00111110011010001000000111010011;
end
if( x <= 32'b10111111100111000010100011110110 && x > 32'b10111111100110101110000101001000)
begin
	y_temp <= 32'b00111110011010100100111100100110;
end
if( x <= 32'b10111111100110101110000101001000 && x > 32'b10111111100110011001100110011010)
begin
	y_temp <= 32'b00111110011011000001111011111100;
end
if( x <= 32'b10111111100110011001100110011010 && x > 32'b10111111100110000101000111101100)
begin
	y_temp <= 32'b00111110011011011111000101010010;
end
if( x <= 32'b10111111100110000101000111101100 && x > 32'b10111111100101110000101000111101)
begin
	y_temp <= 32'b00111110011011111100011000101010;
end
if( x <= 32'b10111111100101110000101000111101 && x > 32'b10111111100101011100001010001111)
begin
	y_temp <= 32'b00111110011100011001110110000010;
end
if( x <= 32'b10111111100101011100001010001111 && x > 32'b10111111100101000111101011100001)
begin
	y_temp <= 32'b00111110011100110111011101011000;
end
if( x <= 32'b10111111100101000111101011100001 && x > 32'b10111111100100110011001100110011)
begin
	y_temp <= 32'b00111110011101010101001110101100;
end
if( x <= 32'b10111111100100110011001100110011 && x > 32'b10111111100100011110101110000101)
begin
	y_temp <= 32'b00111110011101110011001001111101;
end
if( x <= 32'b10111111100100011110101110000101 && x > 32'b10111111100100001010001111010111)
begin
	y_temp <= 32'b00111110011110010001001111001010;
end
if( x <= 32'b10111111100100001010001111010111 && x > 32'b10111111100011110101110000101001)
begin
	y_temp <= 32'b00111110011110101111011110010001;
end
if( x <= 32'b10111111100011110101110000101001 && x > 32'b10111111100011100001010001111011)
begin
	y_temp <= 32'b00111110011111001101110111010001;
end
if( x <= 32'b10111111100011100001010001111011 && x > 32'b10111111100011001100110011001101)
begin
	y_temp <= 32'b00111110011111101100011010001000;
end
if( x <= 32'b10111111100011001100110011001101 && x > 32'b10111111100010111000010100011111)
begin
	y_temp <= 32'b00111110100000000101100011011011;
end
if( x <= 32'b10111111100010111000010100011111 && x > 32'b10111111100010100011110101110001)
begin
	y_temp <= 32'b00111110100000010100111110101100;
end
if( x <= 32'b10111111100010100011110101110001 && x > 32'b10111111100010001111010111000011)
begin
	y_temp <= 32'b00111110100000100100011110110111;
end
if( x <= 32'b10111111100010001111010111000011 && x > 32'b10111111100001111010111000010100)
begin
	y_temp <= 32'b00111110100000110100000011111010;
end
if( x <= 32'b10111111100001111010111000010100 && x > 32'b10111111100001100110011001100110)
begin
	y_temp <= 32'b00111110100001000011101101110101;
end
if( x <= 32'b10111111100001100110011001100110 && x > 32'b10111111100001010001111010111000)
begin
	y_temp <= 32'b00111110100001010011011100100111;
end
if( x <= 32'b10111111100001010001111010111000 && x > 32'b10111111100000111101011100001010)
begin
	y_temp <= 32'b00111110100001100011010000001110;
end
if( x <= 32'b10111111100000111101011100001010 && x > 32'b10111111100000101000111101011100)
begin
	y_temp <= 32'b00111110100001110011001000101010;
end
if( x <= 32'b10111111100000101000111101011100 && x > 32'b10111111100000010100011110101110)
begin
	y_temp <= 32'b00111110100010000011000101111010;
end
if( x <= 32'b10111111100000010100011110101110 && x > 32'b10111111100000000000000000000000)
begin
	y_temp <= 32'b00111110100010010011000111111101;
end
if( x <= 32'b10111111100000000000000000000000 && x > 32'b10111111011111010111000010100100)
begin
	y_temp <= 32'b00111110100010100011001110110001;
end
if( x <= 32'b10111111011111010111000010100100 && x > 32'b10111111011110101110000101001000)
begin
	y_temp <= 32'b00111110100010110011011010010101;
end
if( x <= 32'b10111111011110101110000101001000 && x > 32'b10111111011110000101000111101100)
begin
	y_temp <= 32'b00111110100011000011101010101000;
end
if( x <= 32'b10111111011110000101000111101100 && x > 32'b10111111011101011100001010001111)
begin
	y_temp <= 32'b00111110100011010011111111101001;
end
if( x <= 32'b10111111011101011100001010001111 && x > 32'b10111111011100110011001100110011)
begin
	y_temp <= 32'b00111110100011100100011001010111;
end
if( x <= 32'b10111111011100110011001100110011 && x > 32'b10111111011100001010001111010111)
begin
	y_temp <= 32'b00111110100011110100110111101111;
end
if( x <= 32'b10111111011100001010001111010111 && x > 32'b10111111011011100001010001111011)
begin
	y_temp <= 32'b00111110100100000101011010110010;
end
if( x <= 32'b10111111011011100001010001111011 && x > 32'b10111111011010111000010100011111)
begin
	y_temp <= 32'b00111110100100010110000010011100;
end
if( x <= 32'b10111111011010111000010100011111 && x > 32'b10111111011010001111010111000011)
begin
	y_temp <= 32'b00111110100100100110101110101110;
end
if( x <= 32'b10111111011010001111010111000011 && x > 32'b10111111011001100110011001100110)
begin
	y_temp <= 32'b00111110100100110111011111100100;
end
if( x <= 32'b10111111011001100110011001100110 && x > 32'b10111111011000111101011100001010)
begin
	y_temp <= 32'b00111110100101001000010100111111;
end
if( x <= 32'b10111111011000111101011100001010 && x > 32'b10111111011000010100011110101110)
begin
	y_temp <= 32'b00111110100101011001001110111011;
end
if( x <= 32'b10111111011000010100011110101110 && x > 32'b10111111010111101011100001010010)
begin
	y_temp <= 32'b00111110100101101010001101011000;
end
if( x <= 32'b10111111010111101011100001010010 && x > 32'b10111111010111000010100011110110)
begin
	y_temp <= 32'b00111110100101111011010000010100;
end
if( x <= 32'b10111111010111000010100011110110 && x > 32'b10111111010110011001100110011010)
begin
	y_temp <= 32'b00111110100110001100010111101101;
end
if( x <= 32'b10111111010110011001100110011010 && x > 32'b10111111010101110000101000111101)
begin
	y_temp <= 32'b00111110100110011101100011100001;
end
if( x <= 32'b10111111010101110000101000111101 && x > 32'b10111111010101000111101011100001)
begin
	y_temp <= 32'b00111110100110101110110011101110;
end
if( x <= 32'b10111111010101000111101011100001 && x > 32'b10111111010100011110101110000101)
begin
	y_temp <= 32'b00111110100111000000001000010011;
end
if( x <= 32'b10111111010100011110101110000101 && x > 32'b10111111010011110101110000101001)
begin
	y_temp <= 32'b00111110100111010001100001001110;
end
if( x <= 32'b10111111010011110101110000101001 && x > 32'b10111111010011001100110011001101)
begin
	y_temp <= 32'b00111110100111100010111110011100;
end
if( x <= 32'b10111111010011001100110011001101 && x > 32'b10111111010010100011110101110001)
begin
	y_temp <= 32'b00111110100111110100011111111100;
end
if( x <= 32'b10111111010010100011110101110001 && x > 32'b10111111010001111010111000010100)
begin
	y_temp <= 32'b00111110101000000110000101101100;
end
if( x <= 32'b10111111010001111010111000010100 && x > 32'b10111111010001010001111010111000)
begin
	y_temp <= 32'b00111110101000010111101111101010;
end
if( x <= 32'b10111111010001010001111010111000 && x > 32'b10111111010000101000111101011100)
begin
	y_temp <= 32'b00111110101000101001011101110010;
end
if( x <= 32'b10111111010000101000111101011100 && x > 32'b10111111010000000000000000000000)
begin
	y_temp <= 32'b00111110101000111011010000000101;
end
if( x <= 32'b10111111010000000000000000000000 && x > 32'b10111111001111010111000010100100)
begin
	y_temp <= 32'b00111110101001001101000110011110;
end
if( x <= 32'b10111111001111010111000010100100 && x > 32'b10111111001110101110000101001000)
begin
	y_temp <= 32'b00111110101001011111000000111100;
end
if( x <= 32'b10111111001110101110000101001000 && x > 32'b10111111001110000101000111101100)
begin
	y_temp <= 32'b00111110101001110000111111011101;
end
if( x <= 32'b10111111001110000101000111101100 && x > 32'b10111111001101011100001010001111)
begin
	y_temp <= 32'b00111110101010000011000001111110;
end
if( x <= 32'b10111111001101011100001010001111 && x > 32'b10111111001100110011001100110011)
begin
	y_temp <= 32'b00111110101010010101001000011101;
end
if( x <= 32'b10111111001100110011001100110011 && x > 32'b10111111001100001010001111010111)
begin
	y_temp <= 32'b00111110101010100111010010110111;
end
if( x <= 32'b10111111001100001010001111010111 && x > 32'b10111111001011100001010001111011)
begin
	y_temp <= 32'b00111110101010111001100001001011;
end
if( x <= 32'b10111111001011100001010001111011 && x > 32'b10111111001010111000010100011111)
begin
	y_temp <= 32'b00111110101011001011110011010101;
end
if( x <= 32'b10111111001010111000010100011111 && x > 32'b10111111001010001111010111000011)
begin
	y_temp <= 32'b00111110101011011110001001010011;
end
if( x <= 32'b10111111001010001111010111000011 && x > 32'b10111111001001100110011001100110)
begin
	y_temp <= 32'b00111110101011110000100011000010;
end
if( x <= 32'b10111111001001100110011001100110 && x > 32'b10111111001000111101011100001010)
begin
	y_temp <= 32'b00111110101100000011000000100000;
end
if( x <= 32'b10111111001000111101011100001010 && x > 32'b10111111001000010100011110101110)
begin
	y_temp <= 32'b00111110101100010101100001101010;
end
if( x <= 32'b10111111001000010100011110101110 && x > 32'b10111111000111101011100001010010)
begin
	y_temp <= 32'b00111110101100101000000110011101;
end
if( x <= 32'b10111111000111101011100001010010 && x > 32'b10111111000111000010100011110110)
begin
	y_temp <= 32'b00111110101100111010101110111000;
end
if( x <= 32'b10111111000111000010100011110110 && x > 32'b10111111000110011001100110011010)
begin
	y_temp <= 32'b00111110101101001101011010110110;
end
if( x <= 32'b10111111000110011001100110011010 && x > 32'b10111111000101110000101000111101)
begin
	y_temp <= 32'b00111110101101100000001010010101;
end
if( x <= 32'b10111111000101110000101000111101 && x > 32'b10111111000101000111101011100001)
begin
	y_temp <= 32'b00111110101101110010111101010010;
end
if( x <= 32'b10111111000101000111101011100001 && x > 32'b10111111000100011110101110000101)
begin
	y_temp <= 32'b00111110101110000101110011101011;
end
if( x <= 32'b10111111000100011110101110000101 && x > 32'b10111111000011110101110000101001)
begin
	y_temp <= 32'b00111110101110011000101101011100;
end
if( x <= 32'b10111111000011110101110000101001 && x > 32'b10111111000011001100110011001101)
begin
	y_temp <= 32'b00111110101110101011101010100010;
end
if( x <= 32'b10111111000011001100110011001101 && x > 32'b10111111000010100011110101110001)
begin
	y_temp <= 32'b00111110101110111110101010111011;
end
if( x <= 32'b10111111000010100011110101110001 && x > 32'b10111111000001111010111000010100)
begin
	y_temp <= 32'b00111110101111010001101110100011;
end
if( x <= 32'b10111111000001111010111000010100 && x > 32'b10111111000001010001111010111000)
begin
	y_temp <= 32'b00111110101111100100110101010111;
end
if( x <= 32'b10111111000001010001111010111000 && x > 32'b10111111000000101000111101011100)
begin
	y_temp <= 32'b00111110101111110111111111010101;
end
if( x <= 32'b10111111000000101000111101011100 && x > 32'b10111111000000000000000000000000)
begin
	y_temp <= 32'b00111110110000001011001100011000;
end
if( x <= 32'b10111111000000000000000000000000 && x > 32'b10111110111110101110000101001000)
begin
	y_temp <= 32'b00111110110000011110011100011110;
end
if( x <= 32'b10111110111110101110000101001000 && x > 32'b10111110111101011100001010001111)
begin
	y_temp <= 32'b00111110110000110001101111100011;
end
if( x <= 32'b10111110111101011100001010001111 && x > 32'b10111110111100001010001111010111)
begin
	y_temp <= 32'b00111110110001000101000101100101;
end
if( x <= 32'b10111110111100001010001111010111 && x > 32'b10111110111010111000010100011111)
begin
	y_temp <= 32'b00111110110001011000011110100000;
end
if( x <= 32'b10111110111010111000010100011111 && x > 32'b10111110111001100110011001100110)
begin
	y_temp <= 32'b00111110110001101011111010010000;
end
if( x <= 32'b10111110111001100110011001100110 && x > 32'b10111110111000010100011110101110)
begin
	y_temp <= 32'b00111110110001111111011000110011;
end
if( x <= 32'b10111110111000010100011110101110 && x > 32'b10111110110111000010100011110110)
begin
	y_temp <= 32'b00111110110010010010111010000100;
end
if( x <= 32'b10111110110111000010100011110110 && x > 32'b10111110110101110000101000111101)
begin
	y_temp <= 32'b00111110110010100110011110000001;
end
if( x <= 32'b10111110110101110000101000111101 && x > 32'b10111110110100011110101110000101)
begin
	y_temp <= 32'b00111110110010111010000100100101;
end
if( x <= 32'b10111110110100011110101110000101 && x > 32'b10111110110011001100110011001101)
begin
	y_temp <= 32'b00111110110011001101101101101111;
end
if( x <= 32'b10111110110011001100110011001101 && x > 32'b10111110110001111010111000010100)
begin
	y_temp <= 32'b00111110110011100001011001011000;
end
if( x <= 32'b10111110110001111010111000010100 && x > 32'b10111110110000101000111101011100)
begin
	y_temp <= 32'b00111110110011110101000111100000;
end
if( x <= 32'b10111110110000101000111101011100 && x > 32'b10111110101111010111000010100100)
begin
	y_temp <= 32'b00111110110100001000111000000001;
end
if( x <= 32'b10111110101111010111000010100100 && x > 32'b10111110101110000101000111101100)
begin
	y_temp <= 32'b00111110110100011100101010111000;
end
if( x <= 32'b10111110101110000101000111101100 && x > 32'b10111110101100110011001100110011)
begin
	y_temp <= 32'b00111110110100110000100000000010;
end
if( x <= 32'b10111110101100110011001100110011 && x > 32'b10111110101011100001010001111011)
begin
	y_temp <= 32'b00111110110101000100010111011010;
end
if( x <= 32'b10111110101011100001010001111011 && x > 32'b10111110101010001111010111000011)
begin
	y_temp <= 32'b00111110110101011000010000111110;
end
if( x <= 32'b10111110101010001111010111000011 && x > 32'b10111110101000111101011100001010)
begin
	y_temp <= 32'b00111110110101101100001100101001;
end
if( x <= 32'b10111110101000111101011100001010 && x > 32'b10111110100111101011100001010010)
begin
	y_temp <= 32'b00111110110110000000001010010111;
end
if( x <= 32'b10111110100111101011100001010010 && x > 32'b10111110100110011001100110011010)
begin
	y_temp <= 32'b00111110110110010100001010000110;
end
if( x <= 32'b10111110100110011001100110011010 && x > 32'b10111110100101000111101011100001)
begin
	y_temp <= 32'b00111110110110101000001011110000;
end
if( x <= 32'b10111110100101000111101011100001 && x > 32'b10111110100011110101110000101001)
begin
	y_temp <= 32'b00111110110110111100001111010011;
end
if( x <= 32'b10111110100011110101110000101001 && x > 32'b10111110100010100011110101110001)
begin
	y_temp <= 32'b00111110110111010000010100101010;
end
if( x <= 32'b10111110100010100011110101110001 && x > 32'b10111110100001010001111010111000)
begin
	y_temp <= 32'b00111110110111100100011011110001;
end
if( x <= 32'b10111110100001010001111010111000 && x > 32'b10111110100000000000000000000000)
begin
	y_temp <= 32'b00111110110111111000100100100101;
end
if( x <= 32'b10111110100000000000000000000000 && x > 32'b10111110011101011100001010001111)
begin
	y_temp <= 32'b00111110111000001100101111000010;
end
if( x <= 32'b10111110011101011100001010001111 && x > 32'b10111110011010111000010100011111)
begin
	y_temp <= 32'b00111110111000100000111011000011;
end
if( x <= 32'b10111110011010111000010100011111 && x > 32'b10111110011000010100011110101110)
begin
	y_temp <= 32'b00111110111000110101001000100110;
end
if( x <= 32'b10111110011000010100011110101110 && x > 32'b10111110010101110000101000111101)
begin
	y_temp <= 32'b00111110111001001001010111100101;
end
if( x <= 32'b10111110010101110000101000111101 && x > 32'b10111110010011001100110011001101)
begin
	y_temp <= 32'b00111110111001011101100111111101;
end
if( x <= 32'b10111110010011001100110011001101 && x > 32'b10111110010000101000111101011100)
begin
	y_temp <= 32'b00111110111001110001111001101001;
end
if( x <= 32'b10111110010000101000111101011100 && x > 32'b10111110001110000101000111101100)
begin
	y_temp <= 32'b00111110111010000110001100100111;
end
if( x <= 32'b10111110001110000101000111101100 && x > 32'b10111110001011100001010001111011)
begin
	y_temp <= 32'b00111110111010011010100000110001;
end
if( x <= 32'b10111110001011100001010001111011 && x > 32'b10111110001000111101011100001010)
begin
	y_temp <= 32'b00111110111010101110110110000011;
end
if( x <= 32'b10111110001000111101011100001010 && x > 32'b10111110000110011001100110011010)
begin
	y_temp <= 32'b00111110111011000011001100011011;
end
if( x <= 32'b10111110000110011001100110011010 && x > 32'b10111110000011110101110000101001)
begin
	y_temp <= 32'b00111110111011010111100011110011;
end
if( x <= 32'b10111110000011110101110000101001 && x > 32'b10111110000001010001111010111000)
begin
	y_temp <= 32'b00111110111011101011111100000111;
end
if( x <= 32'b10111110000001010001111010111000 && x > 32'b10111101111101011100001010001111)
begin
	y_temp <= 32'b00111110111100000000010101010011;
end
if( x <= 32'b10111101111101011100001010001111 && x > 32'b10111101111000010100011110101110)
begin
	y_temp <= 32'b00111110111100010100101111010100;
end
if( x <= 32'b10111101111000010100011110101110 && x > 32'b10111101110011001100110011001101)
begin
	y_temp <= 32'b00111110111100101001001010000101;
end
if( x <= 32'b10111101110011001100110011001101 && x > 32'b10111101101110000101000111101100)
begin
	y_temp <= 32'b00111110111100111101100101100001;
end
if( x <= 32'b10111101101110000101000111101100 && x > 32'b10111101101000111101011100001010)
begin
	y_temp <= 32'b00111110111101010010000001100101;
end
if( x <= 32'b10111101101000111101011100001010 && x > 32'b10111101100011110101110000101001)
begin
	y_temp <= 32'b00111110111101100110011110001101;
end
if( x <= 32'b10111101100011110101110000101001 && x > 32'b10111101011101011100001010001111)
begin
	y_temp <= 32'b00111110111101111010111011010100;
end
if( x <= 32'b10111101011101011100001010001111 && x > 32'b10111101010011001100110011001101)
begin
	y_temp <= 32'b00111110111110001111011000110111;
end
if( x <= 32'b10111101010011001100110011001101 && x > 32'b10111101001000111101011100001010)
begin
	y_temp <= 32'b00111110111110100011110110110000;
end
if( x <= 32'b10111101001000111101011100001010 && x > 32'b10111100111101011100001010001111)
begin
	y_temp <= 32'b00111110111110111000010100111101;
end
if( x <= 32'b10111100111101011100001010001111 && x > 32'b10111100101000111101011100001010)
begin
	y_temp <= 32'b00111110111111001100110011011000;
end
if( x <= 32'b10111100101000111101011100001010 && x > 32'b10111100001000111101011100001010)
begin
	y_temp <= 32'b00111110111111100001010001111101;
end
if( x <= 32'b10111100001000111101011100001010 && x > 32'b10101001100011000100111000000000)
begin
	y_temp <= 32'b00111110111111110101110000101001;
end
if( x >= 32'b11000000101000000000000000000000 )
begin
	y_temp <= 0;
end

end
end
assign y = y_temp;

endmodule
